* NGSPICE file created from diff_amp.ext - technology: sky130A

.subckt diff_amp vout gnd vin1 vin2 vdd vinv vamp
X0 Vtail Vtail gnd gnd sky130_fd_pr__nfet_01v8 ad=0.368 pd=2.64 as=0.368 ps=2.64 w=0.92 l=0.16
X1 vs12 vin1 vg34 gnd sky130_fd_pr__nfet_01v8 ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.16
X2 vamp vg34 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.512 pd=3.36 as=0.512 ps=3.36 w=1.28 l=0.16
X3 vamp vin2 vs12 gnd sky130_fd_pr__nfet_01v8 ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.16
X4 vout vinv gnd gnd sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.84 as=0.208 ps=1.84 w=0.52 l=0.16
X5 vout vinv vdd vdd sky130_fd_pr__pfet_01v8 ad=0.416 pd=2.88 as=0.416 ps=2.88 w=1.04 l=0.16
X6 gnd Vtail vs12 gnd sky130_fd_pr__nfet_01v8 ad=0.368 pd=2.64 as=0.368 ps=2.64 w=0.92 l=0.16
X7 vinv vamp vdd vdd sky130_fd_pr__pfet_01v8 ad=0.416 pd=2.88 as=0.416 ps=2.88 w=1.04 l=0.16
X8 vdd vg34 vg34 vdd sky130_fd_pr__pfet_01v8 ad=0.512 pd=3.36 as=0.512 ps=3.36 w=1.28 l=0.16
X9 vinv vamp gnd gnd sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.84 as=0.208 ps=1.84 w=0.52 l=0.16
X10 vdd Vtail gnd sky130_fd_pr__res_xhigh_po w=0.36 l=3
C0 vg34 vin1 0.07432f
C1 vin2 vout 0
C2 vg34 vinv 0
C3 vs12 vin2 0.1312f
C4 vg34 vdd 0.59415f
C5 vout vamp 0
C6 vin2 vamp 0.0921f
C7 Vtail vout 0.02838f
C8 vs12 vamp 0.46352f
C9 Vtail vin2 0.00239f
C10 vin1 vin2 0.02225f
C11 vs12 Vtail 0.05146f
C12 vs12 vin1 0.05358f
C13 vout vinv 0.11673f
C14 vin2 vinv 0
C15 Vtail vamp 0.05528f
C16 vin1 vamp 0
C17 vout vdd 0.38594f
C18 vin2 vdd 0.02223f
C19 vin1 Vtail 0
C20 vs12 vdd 0.00834f
C21 vamp vinv 0.14596f
C22 Vtail vinv 0.03624f
C23 vg34 vout 0
C24 vg34 vin2 0.3161f
C25 vg34 vs12 0.29021f
C26 vamp vdd 0.57504f
C27 Vtail vdd 0.00216f
C28 vin1 vdd 0.00264f
C29 vg34 vamp 0.11337f
C30 vdd vinv 0.52549f
C31 vg34 Vtail 0
C32 vin1 gnd 0.32202f
C33 vin2 gnd 0.32443f
C34 vout gnd 0.26397f
C35 vinv gnd 0.48355f
C36 vamp gnd 0.42931f
C37 vdd gnd 2.29552f
C38 Vtail gnd 1.69512f
C39 vs12 gnd 0.4178f
C40 vg34 gnd 0.51148f
.ends

