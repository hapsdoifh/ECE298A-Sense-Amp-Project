* NGSPICE file created from diff_amp.ext - technology: sky130A

.subckt diff_amp vout gnd vin1 vin2 vdd
X0 Vtail Vtail gnd gnd sky130_fd_pr__nfet_01v8 ad=0.368 pd=2.64 as=0.368 ps=2.64 w=0.92 l=0.16
X1 vs12 vin1 vg34 gnd sky130_fd_pr__nfet_01v8 ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.16
X2 vamp vg34 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.512 pd=3.36 as=0.512 ps=3.36 w=1.28 l=0.16
X3 vamp vin2 vs12 gnd sky130_fd_pr__nfet_01v8 ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.16
X4 vout vinv gnd gnd sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.84 as=0.208 ps=1.84 w=0.52 l=0.16
X5 vout vinv vdd vdd sky130_fd_pr__pfet_01v8 ad=0.416 pd=2.88 as=0.416 ps=2.88 w=1.04 l=0.16
X6 gnd Vtail vs12 gnd sky130_fd_pr__nfet_01v8 ad=0.368 pd=2.64 as=0.368 ps=2.64 w=0.92 l=0.16
X7 vinv vamp vdd vdd sky130_fd_pr__pfet_01v8 ad=0.416 pd=2.88 as=0.416 ps=2.88 w=1.04 l=0.16
X8 vdd vg34 vg34 vdd sky130_fd_pr__pfet_01v8 ad=0.512 pd=3.36 as=0.512 ps=3.36 w=1.28 l=0.16
X9 vinv vamp gnd gnd sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.84 as=0.208 ps=1.84 w=0.52 l=0.16
X10 vdd Vtail gnd sky130_fd_pr__res_xhigh_po w=0.36 l=3
C0 vdd gnd 2.29086f
.ends

