magic
tech sky130A
timestamp 1764392892
<< nwell >>
rect 40 230 150 310
rect -100 -20 690 230
<< nmos >>
rect 370 -150 410 -80
rect 570 -150 610 -80
rect -20 -220 20 -150
rect 170 -220 210 -150
rect 100 -440 140 -370
rect 290 -440 330 -370
<< pmos >>
rect -20 0 20 210
rect 170 0 210 210
rect 370 0 410 210
rect 570 0 610 210
<< ndiff >>
rect 310 -90 370 -80
rect 310 -140 320 -90
rect 340 -140 370 -90
rect 310 -150 370 -140
rect 410 -90 470 -80
rect 410 -140 440 -90
rect 460 -140 470 -90
rect 410 -150 470 -140
rect 510 -90 570 -80
rect 510 -140 520 -90
rect 540 -140 570 -90
rect 510 -150 570 -140
rect 610 -90 670 -80
rect 610 -140 640 -90
rect 660 -140 670 -90
rect 610 -150 670 -140
rect -80 -160 -20 -150
rect -80 -210 -70 -160
rect -50 -210 -20 -160
rect -80 -220 -20 -210
rect 20 -160 80 -150
rect 20 -210 50 -160
rect 70 -210 80 -160
rect 20 -220 80 -210
rect 110 -160 170 -150
rect 110 -210 120 -160
rect 140 -210 170 -160
rect 110 -220 170 -210
rect 210 -160 270 -150
rect 210 -210 240 -160
rect 260 -210 270 -160
rect 210 -220 270 -210
rect 40 -380 100 -370
rect 40 -430 50 -380
rect 70 -430 100 -380
rect 40 -440 100 -430
rect 140 -380 200 -370
rect 140 -430 170 -380
rect 190 -430 200 -380
rect 140 -440 200 -430
rect 230 -380 290 -370
rect 230 -430 240 -380
rect 260 -430 290 -380
rect 230 -440 290 -430
rect 330 -380 390 -370
rect 330 -430 360 -380
rect 380 -430 390 -380
rect 330 -440 390 -430
<< pdiff >>
rect -80 200 -20 210
rect -80 10 -70 200
rect -50 10 -20 200
rect -80 0 -20 10
rect 20 200 80 210
rect 20 10 50 200
rect 70 10 80 200
rect 20 0 80 10
rect 110 200 170 210
rect 110 10 120 200
rect 140 10 170 200
rect 110 0 170 10
rect 210 200 270 210
rect 210 10 240 200
rect 260 10 270 200
rect 210 0 270 10
rect 310 200 370 210
rect 310 10 320 200
rect 340 10 370 200
rect 310 0 370 10
rect 410 200 470 210
rect 410 10 440 200
rect 460 10 470 200
rect 410 0 470 10
rect 510 200 570 210
rect 510 10 520 200
rect 540 10 570 200
rect 510 0 570 10
rect 610 200 670 210
rect 610 10 640 200
rect 660 10 670 200
rect 610 0 670 10
<< ndiffc >>
rect 320 -140 340 -90
rect 440 -140 460 -90
rect 520 -140 540 -90
rect 640 -140 660 -90
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 120 -210 140 -160
rect 240 -210 260 -160
rect 50 -430 70 -380
rect 170 -430 190 -380
rect 240 -430 260 -380
rect 360 -430 380 -380
<< pdiffc >>
rect -70 10 -50 200
rect 50 10 70 200
rect 120 10 140 200
rect 240 10 260 200
rect 320 10 340 200
rect 440 10 460 200
rect 520 10 540 200
rect 640 10 660 200
<< psubdiff >>
rect -90 -400 -30 -380
rect -90 -420 -70 -400
rect -50 -420 -30 -400
rect -90 -440 -30 -420
<< nsubdiff >>
rect 75 275 115 290
rect 75 255 85 275
rect 105 255 115 275
rect 75 240 115 255
<< psubdiffcont >>
rect -70 -420 -50 -400
<< nsubdiffcont >>
rect 85 255 105 275
<< poly >>
rect -20 210 20 240
rect 170 210 210 240
rect 370 210 410 240
rect 570 210 610 240
rect -20 -30 20 0
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 170 -30 210 0
rect 170 -50 180 -30
rect 200 -50 210 -30
rect 170 -60 210 -50
rect 370 -30 410 0
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -80 410 -50
rect 570 -30 610 0
rect 570 -50 580 -30
rect 600 -50 610 -30
rect 570 -80 610 -50
rect 170 -100 210 -90
rect 170 -120 180 -100
rect 200 -120 210 -100
rect -20 -150 20 -130
rect 170 -150 210 -120
rect 370 -170 410 -150
rect 570 -170 610 -150
rect -20 -249 20 -220
rect 170 -240 210 -220
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 100 -320 140 -310
rect 100 -340 110 -320
rect 130 -340 140 -320
rect 100 -370 140 -340
rect 290 -320 330 -310
rect 290 -340 300 -320
rect 320 -340 330 -320
rect 290 -370 330 -340
rect 100 -460 140 -440
rect 290 -460 330 -440
<< polycont >>
rect -10 -50 10 -30
rect 180 -50 200 -30
rect 380 -50 400 -30
rect 580 -50 600 -30
rect 180 -120 200 -100
rect -11 -269 10 -249
rect 110 -340 130 -320
rect 300 -340 320 -320
<< xpolycontact >>
rect 800 90 840 310
rect 730 -310 770 -50
rect 450 -350 670 -310
rect 490 -420 710 -380
rect 510 -520 810 -480
<< xpolyres >>
rect 670 -350 770 -310
rect 800 -380 840 90
rect 450 -480 490 -380
rect 710 -420 840 -380
rect 450 -520 510 -480
<< locali >>
rect 730 300 770 310
rect 75 275 115 285
rect 75 255 85 275
rect 105 255 115 275
rect 75 245 115 255
rect 730 280 740 300
rect 760 280 770 300
rect -80 200 -40 210
rect -80 10 -70 200
rect -50 10 -40 200
rect -80 0 -40 10
rect 40 200 80 210
rect 40 10 50 200
rect 70 10 80 200
rect 40 0 80 10
rect 110 200 150 210
rect 110 10 120 200
rect 140 10 150 200
rect 110 0 150 10
rect 230 200 270 210
rect 230 10 240 200
rect 260 10 270 200
rect 230 0 270 10
rect 310 200 350 210
rect 310 10 320 200
rect 340 10 350 200
rect 310 0 350 10
rect 430 200 470 210
rect 430 10 440 200
rect 460 10 470 200
rect 430 0 470 10
rect 510 200 550 210
rect 510 10 520 200
rect 540 10 550 200
rect 510 0 550 10
rect 630 200 670 210
rect 630 10 640 200
rect 660 10 670 200
rect 730 180 770 280
rect 730 160 740 180
rect 760 160 770 180
rect 730 150 770 160
rect 630 0 670 10
rect -20 -30 20 -20
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 170 -30 210 -20
rect 170 -50 180 -30
rect 200 -50 210 -30
rect 170 -60 210 -50
rect 370 -30 410 -20
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -60 410 -50
rect 570 -30 610 -20
rect 570 -50 580 -30
rect 600 -50 610 -30
rect 570 -60 610 -50
rect 310 -90 350 -80
rect -140 -100 20 -90
rect -140 -120 -130 -100
rect -110 -120 -10 -100
rect 10 -120 20 -100
rect -140 -130 20 -120
rect 170 -100 210 -90
rect 170 -120 180 -100
rect 200 -120 210 -100
rect 170 -130 210 -120
rect 310 -140 320 -90
rect 340 -140 350 -90
rect 310 -150 350 -140
rect 430 -90 470 -80
rect 430 -140 440 -90
rect 460 -140 470 -90
rect 430 -150 470 -140
rect 510 -90 550 -80
rect 510 -140 520 -90
rect 540 -140 550 -90
rect 510 -150 550 -140
rect 630 -90 670 -80
rect 630 -140 640 -90
rect 660 -140 670 -90
rect 630 -150 670 -140
rect -80 -160 -40 -150
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -210 80 -160
rect 40 -220 80 -210
rect 110 -160 150 -150
rect 110 -210 120 -160
rect 140 -210 150 -160
rect 110 -220 150 -210
rect 230 -160 270 -150
rect 230 -210 240 -160
rect 260 -210 270 -160
rect 230 -220 270 -210
rect -20 -249 20 -240
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect -20 -320 140 -310
rect -20 -340 -10 -320
rect 10 -340 110 -320
rect 130 -340 140 -320
rect -20 -350 140 -340
rect 290 -320 330 -310
rect 290 -340 300 -320
rect 320 -340 330 -320
rect 290 -350 330 -340
rect 40 -380 80 -370
rect -90 -400 -30 -380
rect -90 -420 -70 -400
rect -50 -420 -30 -400
rect -90 -440 -30 -420
rect 40 -430 50 -380
rect 70 -430 80 -380
rect 40 -440 80 -430
rect 160 -380 200 -370
rect 160 -430 170 -380
rect 190 -430 200 -380
rect 160 -440 200 -430
rect 230 -380 270 -370
rect 230 -430 240 -380
rect 260 -430 270 -380
rect 230 -440 270 -430
rect 350 -380 390 -370
rect 350 -430 360 -380
rect 380 -430 390 -380
rect 350 -440 390 -430
<< viali >>
rect 85 255 105 275
rect 740 280 760 300
rect -70 10 -50 200
rect 50 10 70 200
rect 120 10 140 200
rect 240 10 260 200
rect 320 10 340 200
rect 440 10 460 200
rect 520 10 540 200
rect 640 10 660 200
rect 740 160 760 180
rect 810 280 830 300
rect -10 -50 10 -30
rect 180 -50 200 -30
rect 380 -50 400 -30
rect 580 -50 600 -30
rect 740 -80 760 -60
rect -130 -120 -110 -100
rect -10 -120 10 -100
rect 180 -120 200 -100
rect 320 -140 340 -90
rect 440 -140 460 -90
rect 520 -140 540 -90
rect 640 -140 660 -90
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 120 -210 140 -160
rect 240 -210 260 -160
rect -11 -269 10 -249
rect -10 -340 10 -320
rect 110 -340 130 -320
rect 300 -340 320 -320
rect 460 -340 480 -320
rect -70 -420 -50 -400
rect 50 -430 70 -380
rect 170 -430 190 -380
rect 240 -430 260 -380
rect 360 -430 380 -380
rect 500 -410 520 -390
rect 600 -510 620 -490
<< metal1 >>
rect -140 300 840 310
rect -140 280 740 300
rect 760 280 810 300
rect 830 280 840 300
rect -140 275 840 280
rect -140 270 85 275
rect 40 255 85 270
rect 105 270 840 275
rect 105 255 150 270
rect 40 230 150 255
rect -80 200 -40 210
rect -80 10 -70 200
rect -50 10 -40 200
rect -80 -20 -40 10
rect 40 200 80 230
rect 40 10 50 200
rect 70 10 80 200
rect 40 0 80 10
rect 110 200 150 230
rect 110 10 120 200
rect 140 10 150 200
rect 110 0 150 10
rect 230 200 270 210
rect 230 10 240 200
rect 260 10 270 200
rect 230 -20 270 10
rect 310 200 350 270
rect 310 10 320 200
rect 340 10 350 200
rect 310 0 350 10
rect 430 200 470 210
rect 430 10 440 200
rect 460 10 470 200
rect -80 -30 210 -20
rect -80 -50 -10 -30
rect 10 -50 180 -30
rect 200 -50 210 -30
rect -80 -60 210 -50
rect 230 -30 410 -20
rect 230 -50 380 -30
rect 400 -50 410 -30
rect 230 -60 410 -50
rect 430 -21 470 10
rect 510 200 550 270
rect 510 10 520 200
rect 540 10 550 200
rect 510 0 550 10
rect 630 210 900 250
rect 630 200 670 210
rect 630 10 640 200
rect 660 10 670 200
rect 510 -21 610 -20
rect 430 -30 610 -21
rect 430 -50 580 -30
rect 600 -50 610 -30
rect 430 -60 610 -50
rect -140 -100 -100 -90
rect -140 -120 -130 -100
rect -110 -120 -100 -100
rect -140 -130 -100 -120
rect -80 -160 -40 -60
rect -20 -100 210 -90
rect -20 -120 -10 -100
rect 10 -120 180 -100
rect 200 -120 210 -100
rect -20 -130 210 -120
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -210 80 -160
rect 40 -220 80 -210
rect 110 -160 150 -150
rect 110 -210 120 -160
rect 140 -210 150 -160
rect 110 -220 150 -210
rect 230 -160 270 -60
rect 230 -210 240 -160
rect 260 -210 270 -160
rect 230 -220 270 -210
rect 310 -90 350 -80
rect 310 -140 320 -90
rect 340 -140 350 -90
rect -140 -249 20 -240
rect -140 -269 -11 -249
rect 10 -269 20 -249
rect -140 -280 20 -269
rect 40 -260 150 -220
rect 310 -250 350 -140
rect 430 -90 470 -60
rect 430 -140 440 -90
rect 460 -140 470 -90
rect 430 -150 470 -140
rect 510 -90 550 -80
rect 510 -140 520 -90
rect 540 -140 550 -90
rect 510 -190 550 -140
rect 630 -90 670 10
rect 730 180 770 190
rect 730 160 740 180
rect 760 160 770 180
rect 730 -60 770 160
rect 730 -80 740 -60
rect 760 -80 770 -60
rect 730 -90 770 -80
rect 630 -140 640 -90
rect 660 -140 670 -90
rect 630 -150 670 -140
rect 510 -230 630 -190
rect -140 -320 20 -310
rect -140 -340 -10 -320
rect 10 -340 20 -320
rect -140 -350 20 -340
rect 40 -380 80 -260
rect 310 -290 570 -250
rect 100 -320 490 -310
rect 100 -340 110 -320
rect 130 -340 300 -320
rect 320 -340 460 -320
rect 480 -340 490 -320
rect 100 -350 490 -340
rect -90 -400 -30 -380
rect -90 -420 -70 -400
rect -50 -420 -30 -400
rect -90 -480 -30 -420
rect 40 -430 50 -380
rect 70 -430 80 -380
rect 40 -440 80 -430
rect 160 -380 200 -370
rect 160 -430 170 -380
rect 190 -430 200 -380
rect 160 -480 200 -430
rect 230 -380 270 -370
rect 230 -430 240 -380
rect 260 -430 270 -380
rect 230 -480 270 -430
rect 350 -380 390 -350
rect 530 -380 570 -290
rect 350 -430 360 -380
rect 380 -430 390 -380
rect 490 -390 570 -380
rect 490 -410 500 -390
rect 520 -410 570 -390
rect 490 -420 570 -410
rect 350 -440 390 -430
rect 590 -480 630 -230
rect -140 -490 630 -480
rect -140 -510 600 -490
rect 620 -510 630 -490
rect -140 -520 630 -510
<< labels >>
rlabel metal1 55 -40 55 -40 1 VG34
rlabel viali -120 -110 -120 -110 1 vin2
rlabel metal1 -61 -261 -57 -255 1 vin1
rlabel metal1 90 -230 90 -230 1 VS12
rlabel metal1 322 -45 334 -35 1 vinv
rlabel metal1 -65 305 -64 306 1 Vdd
rlabel metal1 460 -50 480 -30 1 vinv2
rlabel metal1 320 -190 330 -180 1 vbase
rlabel metal1 90 -520 93 -517 1 Gnd
rlabel metal1 -80 -340 -70 -330 1 vtail
rlabel metal1 870 220 890 240 1 vout
<< end >>
