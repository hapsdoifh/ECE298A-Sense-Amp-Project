magic
tech sky130A
timestamp 1762137474
<< error_p >>
rect -18 62 18 72
rect -36 54 -28 62
rect -26 54 26 62
rect 28 54 36 62
rect -44 50 -10 54
rect -44 46 -32 50
rect -18 46 -10 50
rect 10 50 44 54
rect 10 46 18 50
rect 32 46 44 50
rect -36 -46 -32 46
rect 32 -46 36 46
rect -73 -54 -65 -46
rect -59 -54 -51 -46
rect -44 -49 -32 -46
rect -18 -49 -10 -46
rect 10 -49 18 -46
rect 32 -49 44 -46
rect -44 -54 44 -49
rect -81 -56 -43 -54
rect -36 -56 -28 -54
rect -26 -56 26 -54
rect -81 -59 26 -56
rect -81 -62 -43 -59
rect -36 -62 -28 -59
rect -26 -62 26 -59
rect 28 -62 36 -54
rect -73 -68 -51 -62
rect -18 -68 18 -62
rect -81 -76 -43 -68
rect -36 -76 -28 -68
rect -26 -72 26 -68
rect -26 -76 -18 -72
rect 18 -76 26 -72
rect 28 -76 36 -68
rect -73 -84 -65 -76
rect -59 -84 -51 -76
rect -44 -80 -10 -76
rect -44 -84 -32 -80
rect -18 -84 -10 -80
rect 10 -80 44 -76
rect 10 -84 18 -80
rect 32 -84 44 -80
rect -36 -116 -32 -84
rect 32 -116 36 -84
rect -44 -120 -32 -116
rect -18 -120 -10 -116
rect -44 -124 -10 -120
rect 10 -120 18 -116
rect 32 -120 44 -116
rect 10 -124 44 -120
rect -36 -132 -28 -124
rect -26 -132 -18 -124
rect 18 -132 26 -124
rect 28 -132 36 -124
rect -10 -137 9 -136
<< nmos >>
rect -10 -124 9 -76
<< pmos >>
rect -10 -54 9 54
<< ndiff >>
rect -18 -124 -10 -76
rect 9 -124 18 -76
<< pdiff >>
rect -18 -54 -10 54
rect 9 -54 18 54
<< ndiffc >>
rect -36 -124 -18 -76
rect 18 -124 36 -76
<< pdiffc >>
rect -36 -54 -18 54
rect 18 -54 36 54
<< poly >>
rect -10 54 9 66
rect -10 -59 9 -54
rect -51 -71 9 -59
rect -10 -76 9 -71
rect -10 -136 9 -124
<< polycont >>
rect -73 -76 -51 -54
<< metal1 >>
rect -54 72 54 104
rect -36 54 -18 72
<< end >>
