* SPICE3 file created from diff_amp.ext - technology: sky130A

X0 Gnd vtail VS12 Gnd sky130_fd_pr__nfet_01v8 ad=0.54 pd=3 as=0.54 ps=3 w=0.9 l=0.4
X1 vout vinv2 Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.2 as=0.3 ps=2.2 w=0.5 l=0.4
X2 VS12 vin1 VG34 Gnd sky130_fd_pr__nfet_01v8 ad=1.08 pd=4.8 as=1.08 ps=4.8 w=1.8 l=0.4
X3 vinv2 vinv Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.2 as=0.6 ps=3.2 w=1 l=0.4
X4 Vdd VG34 VG34 Vdd sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.4 as=0.36 ps=2.4 w=0.6 l=0.4
X5 vtail vtail Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.54 pd=3 as=0.54 ps=3 w=0.9 l=0.4
X6 vout vinv2 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.2 as=0.6 ps=3.2 w=1 l=0.4
X7 vinv vin2 VS12 Gnd sky130_fd_pr__nfet_01v8 ad=1.08 pd=4.8 as=1.08 ps=4.8 w=1.8 l=0.4
X8 vinv VG34 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.4 as=0.36 ps=2.4 w=0.6 l=0.4
X9 vinv2 vinv Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.2 as=0.3 ps=2.2 w=0.5 l=0.4
X10 Vdd vtail Gnd sky130_fd_pr__res_xhigh_po w=0.4 l=0.96
C0 Vdd Gnd 2.22558f 
