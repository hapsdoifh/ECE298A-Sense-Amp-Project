magic
tech sky130A
timestamp 1763530409
<< nwell >>
rect -100 -20 380 160
<< nmos >>
rect -20 -220 20 -150
rect 260 -220 300 -150
rect 180 -440 220 -370
<< pmos >>
rect -20 0 20 140
rect 260 0 300 140
<< ndiff >>
rect -80 -160 -20 -150
rect -80 -210 -70 -160
rect -50 -210 -20 -160
rect -80 -220 -20 -210
rect 20 -160 80 -150
rect 20 -210 50 -160
rect 70 -210 80 -160
rect 20 -220 80 -210
rect 200 -160 260 -150
rect 200 -210 210 -160
rect 230 -210 260 -160
rect 200 -220 260 -210
rect 300 -160 360 -150
rect 300 -210 330 -160
rect 350 -210 360 -160
rect 300 -220 360 -210
rect 120 -380 180 -370
rect 120 -430 130 -380
rect 150 -430 180 -380
rect 120 -440 180 -430
rect 220 -380 280 -370
rect 220 -430 250 -380
rect 270 -430 280 -380
rect 220 -440 280 -430
<< pdiff >>
rect -80 130 -20 140
rect -80 10 -70 130
rect -50 10 -20 130
rect -80 0 -20 10
rect 20 130 80 140
rect 20 10 50 130
rect 70 10 80 130
rect 200 130 260 140
rect 20 0 80 10
rect 200 10 210 130
rect 230 10 260 130
rect 200 0 260 10
rect 300 130 360 140
rect 300 10 330 130
rect 350 10 360 130
rect 300 0 360 10
<< ndiffc >>
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 210 -210 230 -160
rect 330 -210 350 -160
rect 130 -430 150 -380
rect 250 -430 270 -380
<< pdiffc >>
rect -70 10 -50 130
rect 50 10 70 130
rect 210 10 230 130
rect 330 10 350 130
<< psubdiff >>
rect 0 -350 80 -330
rect 0 -390 20 -350
rect 60 -390 80 -350
rect 0 -410 80 -390
<< nsubdiff >>
rect 115 90 165 105
rect 115 70 130 90
rect 150 70 165 90
rect 115 55 165 70
<< psubdiffcont >>
rect 20 -390 60 -350
<< nsubdiffcont >>
rect 130 70 150 90
<< poly >>
rect -20 140 20 170
rect 260 140 300 170
rect -20 -30 20 0
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 260 -30 300 0
rect 260 -50 270 -30
rect 290 -50 300 -30
rect 260 -60 300 -50
rect -20 -100 20 -90
rect -20 -120 -10 -100
rect 10 -120 20 -100
rect -20 -150 20 -120
rect 260 -150 300 -130
rect -20 -240 20 -220
rect 260 -249 300 -220
rect 260 -269 269 -249
rect 290 -269 300 -249
rect 260 -280 300 -269
rect 180 -320 220 -310
rect 180 -340 190 -320
rect 210 -340 220 -320
rect 180 -370 220 -340
rect 180 -460 220 -440
<< polycont >>
rect -10 -50 10 -30
rect 270 -50 290 -30
rect -10 -120 10 -100
rect 269 -269 290 -249
rect 190 -340 210 -320
<< locali >>
rect -80 130 -40 140
rect -80 10 -71 130
rect -50 10 -40 130
rect -80 0 -40 10
rect 40 130 80 140
rect 40 10 50 130
rect 70 10 80 130
rect 200 130 240 140
rect 120 90 160 100
rect 120 70 130 90
rect 150 70 160 90
rect 120 60 160 70
rect 40 0 80 10
rect 200 10 210 130
rect 230 10 240 130
rect 200 0 240 10
rect 320 130 360 140
rect 320 10 330 130
rect 350 10 360 130
rect 320 0 360 10
rect -20 -30 20 -20
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 260 -30 300 -20
rect 260 -50 270 -30
rect 290 -50 300 -30
rect 260 -60 300 -50
rect -20 -100 20 -90
rect -20 -120 -10 -100
rect 10 -120 20 -100
rect -20 -130 20 -120
rect 260 -100 420 -90
rect 260 -120 270 -100
rect 290 -120 390 -100
rect 410 -120 420 -100
rect 260 -130 420 -120
rect -80 -160 -40 -150
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -210 80 -160
rect 40 -220 80 -210
rect 200 -160 240 -150
rect 200 -210 210 -160
rect 230 -210 240 -160
rect 200 -220 240 -210
rect 320 -160 360 -150
rect 320 -210 330 -160
rect 350 -210 360 -160
rect 320 -220 360 -210
rect 260 -249 300 -240
rect 260 -269 269 -249
rect 290 -269 300 -249
rect 260 -280 300 -269
rect 180 -320 220 -310
rect 0 -350 80 -330
rect 180 -340 190 -320
rect 210 -340 220 -320
rect 180 -350 220 -340
rect 0 -390 20 -350
rect 60 -390 80 -350
rect 0 -410 80 -390
rect 120 -380 160 -370
rect 120 -430 130 -380
rect 150 -430 160 -380
rect 120 -440 160 -430
rect 240 -380 280 -370
rect 240 -430 250 -380
rect 270 -430 280 -380
rect 240 -440 280 -430
<< viali >>
rect -71 10 -70 130
rect -70 10 -50 130
rect 50 10 70 130
rect 130 70 150 90
rect 210 10 230 130
rect 330 10 350 130
rect -10 -50 10 -30
rect 270 -50 290 -30
rect -10 -120 10 -100
rect 270 -120 290 -100
rect 390 -120 410 -100
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 210 -210 230 -160
rect 330 -210 350 -160
rect 269 -269 290 -249
rect 190 -340 210 -320
rect 20 -390 60 -350
rect 130 -430 150 -380
rect 250 -430 270 -380
<< metal1 >>
rect -100 200 380 270
rect -80 130 -40 140
rect -80 10 -71 130
rect -50 10 -40 130
rect -80 -20 -40 10
rect 40 130 80 200
rect 40 10 50 130
rect 70 10 80 130
rect 120 90 160 200
rect 120 70 130 90
rect 150 70 160 90
rect 120 60 160 70
rect 200 130 240 200
rect 40 0 80 10
rect 200 10 210 130
rect 230 10 240 130
rect 200 0 240 10
rect 320 130 360 140
rect 320 10 330 130
rect 350 10 360 130
rect 320 -20 360 10
rect -80 -30 300 -20
rect -80 -50 -10 -30
rect 10 -50 270 -30
rect 290 -50 300 -30
rect -80 -60 300 -50
rect 320 -60 420 -20
rect -80 -160 -40 -60
rect -20 -100 300 -90
rect -20 -120 -10 -100
rect 10 -120 270 -100
rect 290 -120 300 -100
rect -20 -130 300 -120
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -210 80 -160
rect 40 -240 80 -210
rect 200 -160 240 -150
rect 200 -210 210 -160
rect 230 -210 240 -160
rect 200 -240 240 -210
rect 320 -160 360 -60
rect 380 -100 420 -90
rect 380 -120 390 -100
rect 410 -120 420 -100
rect 380 -130 420 -120
rect 320 -210 330 -160
rect 350 -210 360 -160
rect 320 -220 360 -210
rect 40 -280 240 -240
rect 260 -249 420 -240
rect 260 -269 269 -249
rect 290 -269 420 -249
rect 260 -280 420 -269
rect 0 -350 80 -330
rect 0 -390 20 -350
rect 60 -390 80 -350
rect 0 -470 80 -390
rect 120 -380 160 -280
rect 180 -320 420 -310
rect 180 -340 190 -320
rect 210 -340 420 -320
rect 180 -350 420 -340
rect 120 -430 130 -380
rect 150 -430 160 -380
rect 120 -440 160 -430
rect 240 -380 280 -370
rect 240 -430 250 -380
rect 270 -430 280 -380
rect 240 -470 280 -430
rect -100 -540 380 -470
<< labels >>
rlabel metal1 55 -40 55 -40 1 VG34
rlabel metal1 341 -76 341 -76 1 Vout
rlabel metal1 90 -510 93 -507 1 Gnd
rlabel metal1 340 -260 340 -260 1 Vin2
rlabel viali 400 -110 400 -110 1 vin1
rlabel metal1 -65 235 -64 236 1 Vdd
rlabel metal1 370 -330 370 -330 1 Vtail
<< end >>
