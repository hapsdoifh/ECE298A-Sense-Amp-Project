magic
tech sky130A
timestamp 1764201597
<< nwell >>
rect 40 160 150 240
rect -100 -20 690 160
<< nmos >>
rect 370 -150 410 -80
rect 570 -150 610 -80
rect -20 -220 20 -150
rect 170 -220 210 -150
rect 60 -350 130 -310
<< pmos >>
rect -20 0 20 140
rect 170 0 210 140
rect 370 0 410 140
rect 570 0 610 140
<< ndiff >>
rect 310 -90 370 -80
rect 310 -140 320 -90
rect 340 -140 370 -90
rect 310 -150 370 -140
rect 410 -90 470 -80
rect 410 -140 440 -90
rect 460 -140 470 -90
rect 410 -150 470 -140
rect 510 -90 570 -80
rect 510 -140 520 -90
rect 540 -140 570 -90
rect 510 -150 570 -140
rect 610 -90 670 -80
rect 610 -140 640 -90
rect 660 -140 670 -90
rect 610 -150 670 -140
rect -80 -160 -20 -150
rect -80 -210 -70 -160
rect -50 -210 -20 -160
rect -80 -220 -20 -210
rect 20 -160 80 -150
rect 20 -210 50 -160
rect 70 -210 80 -160
rect 20 -220 80 -210
rect 110 -160 170 -150
rect 110 -210 120 -160
rect 140 -210 170 -160
rect 110 -220 170 -210
rect 210 -160 270 -150
rect 210 -210 240 -160
rect 260 -210 270 -160
rect 210 -220 270 -210
rect 60 -260 130 -250
rect 60 -280 70 -260
rect 120 -280 130 -260
rect 60 -310 130 -280
rect 60 -380 130 -350
rect 60 -400 70 -380
rect 120 -400 130 -380
rect 60 -410 130 -400
<< pdiff >>
rect -80 130 -20 140
rect -80 10 -70 130
rect -50 10 -20 130
rect -80 0 -20 10
rect 20 130 80 140
rect 20 10 50 130
rect 70 10 80 130
rect 20 0 80 10
rect 110 130 170 140
rect 110 10 120 130
rect 140 10 170 130
rect 110 0 170 10
rect 210 130 270 140
rect 210 10 240 130
rect 260 10 270 130
rect 210 0 270 10
rect 310 130 370 140
rect 310 10 320 130
rect 340 10 370 130
rect 310 0 370 10
rect 410 130 470 140
rect 410 10 440 130
rect 460 10 470 130
rect 410 0 470 10
rect 510 130 570 140
rect 510 10 520 130
rect 540 10 570 130
rect 510 0 570 10
rect 610 130 670 140
rect 610 10 640 130
rect 660 10 670 130
rect 610 0 670 10
<< ndiffc >>
rect 320 -140 340 -90
rect 440 -140 460 -90
rect 520 -140 540 -90
rect 640 -140 660 -90
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 120 -210 140 -160
rect 240 -210 260 -160
rect 70 -280 120 -260
rect 70 -400 120 -380
<< pdiffc >>
rect -70 10 -50 130
rect 50 10 70 130
rect 120 10 140 130
rect 240 10 260 130
rect 320 10 340 130
rect 440 10 460 130
rect 520 10 540 130
rect 640 10 660 130
<< psubdiff >>
rect 180 -330 240 -310
rect 180 -350 200 -330
rect 220 -350 240 -330
rect 180 -370 240 -350
<< nsubdiff >>
rect 75 205 115 220
rect 75 185 85 205
rect 105 185 115 205
rect 75 170 115 185
<< psubdiffcont >>
rect 200 -350 220 -330
<< nsubdiffcont >>
rect 85 185 105 205
<< poly >>
rect -20 140 20 170
rect 170 140 210 170
rect 370 140 410 170
rect 570 140 610 170
rect -20 -30 20 0
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 170 -30 210 0
rect 170 -50 180 -30
rect 200 -50 210 -30
rect 170 -60 210 -50
rect 370 -30 410 0
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -80 410 -50
rect 570 -30 610 0
rect 570 -50 580 -30
rect 600 -50 610 -30
rect 570 -80 610 -50
rect 170 -100 210 -90
rect 170 -120 180 -100
rect 200 -120 210 -100
rect -20 -150 20 -130
rect 170 -150 210 -120
rect 370 -170 410 -150
rect 570 -170 610 -150
rect -20 -249 20 -220
rect 170 -240 210 -220
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 0 -320 60 -310
rect 0 -340 10 -320
rect 30 -340 60 -320
rect 0 -350 60 -340
rect 130 -350 150 -310
<< polycont >>
rect -10 -50 10 -30
rect 180 -50 200 -30
rect 380 -50 400 -30
rect 580 -50 600 -30
rect 180 -120 200 -100
rect -11 -269 10 -249
rect 10 -340 30 -320
<< locali >>
rect 75 205 115 215
rect 75 185 85 205
rect 105 185 115 205
rect 75 175 115 185
rect -80 130 -40 140
rect -80 10 -70 130
rect -50 10 -40 130
rect -80 0 -40 10
rect 40 130 80 140
rect 40 10 50 130
rect 70 10 80 130
rect 40 0 80 10
rect 110 130 150 140
rect 110 10 120 130
rect 140 10 150 130
rect 110 0 150 10
rect 230 130 270 140
rect 230 10 240 130
rect 260 10 270 130
rect 230 0 270 10
rect 310 130 350 140
rect 310 10 320 130
rect 340 10 350 130
rect 310 0 350 10
rect 430 130 470 140
rect 430 10 440 130
rect 460 10 470 130
rect 430 0 470 10
rect 510 130 550 140
rect 510 10 520 130
rect 540 10 550 130
rect 510 0 550 10
rect 630 130 670 140
rect 630 10 640 130
rect 660 10 670 130
rect 630 0 670 10
rect -20 -30 20 -20
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 170 -30 210 -20
rect 170 -50 180 -30
rect 200 -50 210 -30
rect 170 -60 210 -50
rect 370 -30 410 -20
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -60 410 -50
rect 570 -30 610 -20
rect 570 -50 580 -30
rect 600 -50 610 -30
rect 570 -60 610 -50
rect 310 -90 350 -80
rect -140 -100 20 -90
rect -140 -120 -130 -100
rect -110 -120 -10 -100
rect 10 -120 20 -100
rect -140 -130 20 -120
rect 170 -100 210 -90
rect 170 -120 180 -100
rect 200 -120 210 -100
rect 170 -130 210 -120
rect 310 -140 320 -90
rect 340 -140 350 -90
rect 310 -150 350 -140
rect 430 -90 470 -80
rect 430 -140 440 -90
rect 460 -140 470 -90
rect 430 -150 470 -140
rect 510 -90 550 -80
rect 510 -140 520 -90
rect 540 -140 550 -90
rect 510 -150 550 -140
rect 630 -90 670 -80
rect 630 -140 640 -90
rect 660 -140 670 -90
rect 630 -150 670 -140
rect -80 -160 -40 -150
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -210 80 -160
rect 40 -220 80 -210
rect 110 -160 150 -150
rect 110 -210 120 -160
rect 140 -210 150 -160
rect 110 -220 150 -210
rect 230 -160 270 -150
rect 230 -210 240 -160
rect 260 -210 270 -160
rect 230 -220 270 -210
rect -20 -249 20 -240
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 60 -260 130 -250
rect 60 -280 70 -260
rect 120 -280 130 -260
rect 60 -290 130 -280
rect 310 -280 470 -270
rect 310 -300 320 -280
rect 340 -300 440 -280
rect 460 -300 470 -280
rect 310 -310 470 -300
rect 0 -320 40 -310
rect 0 -340 10 -320
rect 30 -340 40 -320
rect 0 -350 40 -340
rect 180 -330 240 -310
rect 180 -350 200 -330
rect 220 -350 240 -330
rect 180 -370 240 -350
rect 60 -380 130 -370
rect 60 -400 70 -380
rect 120 -400 130 -380
rect 60 -410 130 -400
<< viali >>
rect 85 185 105 205
rect -70 10 -50 130
rect 50 10 70 130
rect 120 10 140 130
rect 240 10 260 130
rect 320 10 340 130
rect 440 10 460 130
rect 520 10 540 130
rect 640 10 660 130
rect -10 -50 10 -30
rect 180 -50 200 -30
rect 380 -50 400 -30
rect 580 -50 600 -30
rect -130 -120 -110 -100
rect -10 -120 10 -100
rect 180 -120 200 -100
rect 320 -140 340 -90
rect 440 -140 460 -90
rect 520 -140 540 -90
rect 640 -140 660 -90
rect -70 -210 -50 -160
rect 50 -210 70 -160
rect 120 -210 140 -160
rect 240 -210 260 -160
rect -11 -269 10 -249
rect 70 -280 120 -260
rect 320 -300 340 -280
rect 440 -300 460 -280
rect 10 -340 30 -320
rect 200 -350 220 -330
rect 70 -400 120 -380
<< metal1 >>
rect -140 205 670 240
rect -140 200 85 205
rect 40 185 85 200
rect 105 200 670 205
rect 105 185 150 200
rect 40 160 150 185
rect -80 130 -40 140
rect -80 10 -70 130
rect -50 10 -40 130
rect -80 -20 -40 10
rect 40 130 80 160
rect 40 10 50 130
rect 70 10 80 130
rect 40 0 80 10
rect 110 130 150 160
rect 110 10 120 130
rect 140 10 150 130
rect 110 0 150 10
rect 230 130 270 140
rect 230 10 240 130
rect 260 10 270 130
rect 230 -20 270 10
rect 310 130 350 200
rect 310 10 320 130
rect 340 10 350 130
rect 310 0 350 10
rect 430 130 470 140
rect 430 10 440 130
rect 460 10 470 130
rect -80 -30 210 -20
rect -80 -50 -10 -30
rect 10 -50 180 -30
rect 200 -50 210 -30
rect -80 -60 210 -50
rect 230 -30 410 -20
rect 230 -50 380 -30
rect 400 -50 410 -30
rect 230 -60 410 -50
rect 430 -21 470 10
rect 510 130 550 200
rect 510 10 520 130
rect 540 10 550 130
rect 510 0 550 10
rect 630 130 670 140
rect 630 10 640 130
rect 660 10 670 130
rect 510 -21 610 -20
rect 430 -30 610 -21
rect 430 -50 580 -30
rect 600 -50 610 -30
rect 430 -60 610 -50
rect -140 -100 -100 -90
rect -140 -120 -130 -100
rect -110 -120 -100 -100
rect -140 -130 -100 -120
rect -80 -160 -40 -60
rect -20 -100 210 -90
rect -20 -120 -10 -100
rect 10 -120 180 -100
rect 200 -120 210 -100
rect -20 -130 210 -120
rect -80 -210 -70 -160
rect -50 -210 -40 -160
rect -80 -220 -40 -210
rect 40 -160 80 -150
rect 40 -210 50 -160
rect 70 -210 80 -160
rect 40 -220 80 -210
rect 110 -160 150 -150
rect 110 -210 120 -160
rect 140 -210 150 -160
rect 110 -220 150 -210
rect 230 -160 270 -60
rect 230 -210 240 -160
rect 260 -210 270 -160
rect 230 -220 270 -210
rect 310 -90 350 -80
rect 310 -140 320 -90
rect 340 -140 350 -90
rect -140 -249 20 -240
rect -140 -269 -11 -249
rect 10 -269 20 -249
rect 40 -250 150 -220
rect -140 -280 20 -269
rect 60 -260 130 -250
rect 60 -280 70 -260
rect 120 -280 130 -260
rect 60 -290 130 -280
rect 310 -280 350 -140
rect 430 -90 470 -60
rect 430 -140 440 -90
rect 460 -140 470 -90
rect 430 -150 470 -140
rect 510 -90 550 -80
rect 510 -140 520 -90
rect 540 -140 550 -90
rect 510 -190 550 -140
rect 630 -90 670 10
rect 630 -140 640 -90
rect 660 -140 670 -90
rect 630 -150 670 -140
rect 310 -300 320 -280
rect 340 -300 350 -280
rect 310 -310 350 -300
rect 370 -230 550 -190
rect -140 -320 40 -310
rect -140 -340 10 -320
rect 30 -340 40 -320
rect -140 -350 40 -340
rect 180 -330 240 -310
rect 370 -330 410 -230
rect 430 -280 470 -270
rect 430 -300 440 -280
rect 460 -300 470 -280
rect 430 -310 470 -300
rect 180 -350 200 -330
rect 220 -350 410 -330
rect 180 -370 410 -350
rect 60 -380 130 -370
rect 60 -400 70 -380
rect 120 -400 130 -380
rect 60 -410 130 -400
rect 180 -410 240 -370
rect -140 -450 240 -410
<< labels >>
rlabel metal1 55 -40 55 -40 1 VG34
rlabel viali -120 -110 -120 -110 1 vin2
rlabel metal1 -61 -261 -57 -255 1 vin1
rlabel metal1 90 -450 93 -447 1 Gnd
rlabel metal1 90 -230 90 -230 1 VS12
rlabel metal1 -30 -330 -30 -330 1 Vtail
rlabel metal1 470 -50 480 -40 1 Vout2
rlabel metal1 322 -45 334 -35 1 vinv
rlabel metal1 320 -250 340 -230 1 vbase
rlabel metal1 650 -51 660 -40 1 voutf
rlabel metal1 -65 235 -64 236 1 Vdd
<< end >>
