* SPICE3 file created from diff_amp.ext - technology: sky130A

X0 VS12 vin1 VG34 Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X1 vinv VG34 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=5.4 as=1.26 ps=5.4 w=2.1 l=0.4
X2 voutf Vout2 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=5.4 as=1.26 ps=5.4 w=2.1 l=0.4
X3 Vdd vbase Gnd sky130_fd_pr__res_xhigh_po w=0.4 l=7.96
X4 VS12 Vtail Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X5 Vdd VG34 VG34 Vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=5.4 as=1.26 ps=5.4 w=2.1 l=0.4
X6 vbase Gnd Gnd sky130_fd_pr__res_xhigh_po w=0.4 l=1.56
X7 Vout2 vinv vbase Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X8 voutf Vout2 Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X9 vinv vin2 VS12 Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X10 Vout2 vinv Vdd Vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=5.4 as=1.26 ps=5.4 w=2.1 l=0.4
C0 Vdd Gnd 3.33134f
