magic
tech sky130A
timestamp 1764725471
<< nwell >>
rect -4 312 96 332
rect -4 304 452 312
rect -48 268 452 304
rect -100 124 452 268
rect -100 100 168 124
rect -100 76 136 100
<< nmos >>
rect 216 12 232 64
rect 340 12 356 64
rect -32 -204 -16 -24
rect 92 -204 108 -24
rect 216 -204 232 -112
rect 340 -204 356 -112
<< pmos >>
rect -32 120 -16 248
rect 92 120 108 248
rect 216 144 232 248
rect 340 144 356 248
<< ndiff >>
rect 176 56 216 64
rect 176 20 184 56
rect 204 20 216 56
rect 176 12 216 20
rect 232 56 272 64
rect 232 20 244 56
rect 264 20 272 56
rect 232 12 272 20
rect 300 56 340 64
rect 300 20 308 56
rect 328 20 340 56
rect 300 12 340 20
rect 356 56 396 64
rect 356 20 368 56
rect 388 20 396 56
rect 356 12 396 20
rect -72 -32 -32 -24
rect -72 -196 -64 -32
rect -44 -196 -32 -32
rect -72 -204 -32 -196
rect -16 -32 24 -24
rect -16 -196 -4 -32
rect 16 -196 24 -32
rect -16 -204 24 -196
rect 52 -32 92 -24
rect 52 -196 60 -32
rect 80 -196 92 -32
rect 52 -204 92 -196
rect 108 -32 148 -24
rect 108 -196 120 -32
rect 140 -196 148 -32
rect 108 -204 148 -196
rect 176 -120 216 -112
rect 176 -196 184 -120
rect 204 -196 216 -120
rect 176 -204 216 -196
rect 232 -120 272 -112
rect 232 -196 244 -120
rect 264 -196 272 -120
rect 232 -204 272 -196
rect 300 -120 340 -112
rect 300 -196 308 -120
rect 328 -196 340 -120
rect 300 -204 340 -196
rect 356 -120 396 -112
rect 356 -196 368 -120
rect 388 -196 396 -120
rect 356 -204 396 -196
<< pdiff >>
rect -72 240 -32 248
rect -72 128 -64 240
rect -44 128 -32 240
rect -72 120 -32 128
rect -16 240 24 248
rect -16 128 -4 240
rect 16 128 24 240
rect -16 120 24 128
rect 52 240 92 248
rect 52 128 60 240
rect 80 128 92 240
rect 52 120 92 128
rect 108 240 148 248
rect 108 128 120 240
rect 140 128 148 240
rect 176 240 216 248
rect 176 152 184 240
rect 204 152 216 240
rect 176 144 216 152
rect 232 240 272 248
rect 232 152 244 240
rect 264 152 272 240
rect 232 144 272 152
rect 300 240 340 248
rect 300 152 308 240
rect 328 152 340 240
rect 300 144 340 152
rect 356 240 396 248
rect 356 152 368 240
rect 388 152 396 240
rect 356 144 396 152
rect 108 120 148 128
<< ndiffc >>
rect 184 20 204 56
rect 244 20 264 56
rect 308 20 328 56
rect 368 20 388 56
rect -64 -196 -44 -32
rect -4 -196 16 -32
rect 60 -196 80 -32
rect 120 -196 140 -32
rect 184 -196 204 -120
rect 244 -196 264 -120
rect 308 -196 328 -120
rect 368 -196 388 -120
<< pdiffc >>
rect -64 128 -44 240
rect -4 128 16 240
rect 60 128 80 240
rect 120 128 140 240
rect 184 152 204 240
rect 244 152 264 240
rect 308 152 328 240
rect 368 152 388 240
<< psubdiff >>
rect -88 -320 -28 -300
rect -88 -340 -68 -320
rect -48 -340 -28 -320
rect -88 -360 -28 -340
<< nsubdiff >>
rect 24 304 68 312
rect 24 284 36 304
rect 56 284 68 304
rect 24 276 68 284
<< psubdiffcont >>
rect -68 -340 -48 -320
<< nsubdiffcont >>
rect 36 284 56 304
<< poly >>
rect -32 248 -16 264
rect 92 248 108 264
rect 216 248 232 264
rect 340 248 356 264
rect 216 124 232 144
rect 340 124 356 144
rect -32 100 -16 120
rect 92 100 108 120
rect 204 116 244 124
rect -44 92 -4 100
rect -44 68 -36 92
rect -12 68 -4 92
rect -44 60 -4 68
rect 80 92 120 100
rect 80 68 88 92
rect 112 68 120 92
rect 204 92 212 116
rect 236 92 244 116
rect 204 84 244 92
rect 328 116 368 124
rect 328 92 336 116
rect 360 92 368 116
rect 328 84 368 92
rect 80 60 120 68
rect 216 64 232 84
rect 340 64 356 84
rect 80 28 120 36
rect 80 4 88 28
rect 112 4 120 28
rect 80 -4 120 4
rect -32 -24 -16 -4
rect 92 -24 108 -4
rect 216 -8 232 12
rect 340 -8 356 12
rect 204 -60 244 -52
rect 204 -84 212 -60
rect 236 -84 244 -60
rect 204 -92 244 -84
rect 328 -60 368 -52
rect 328 -84 336 -60
rect 360 -84 368 -60
rect 328 -92 368 -84
rect 216 -112 232 -92
rect 340 -112 356 -92
rect -32 -224 -16 -204
rect 92 -224 108 -204
rect 216 -220 232 -204
rect 340 -220 356 -204
rect -44 -232 -4 -224
rect -44 -256 -36 -232
rect -12 -256 -4 -232
rect -44 -264 -4 -256
<< polycont >>
rect -36 68 -12 92
rect 88 68 112 92
rect 212 92 236 116
rect 336 92 360 116
rect 88 4 112 28
rect 212 -84 236 -60
rect 336 -84 360 -60
rect -36 -256 -12 -232
<< xpolycontact >>
rect 452 -20 488 320
rect 148 -304 452 -268
<< xpolyres >>
rect 452 -304 488 -20
<< locali >>
rect 28 304 64 312
rect 28 284 36 304
rect 56 284 64 304
rect 28 276 64 284
rect -72 240 -36 248
rect -72 128 -64 240
rect -44 128 -36 240
rect -72 120 -36 128
rect -12 240 24 248
rect -12 128 -4 240
rect 16 128 24 240
rect -12 120 24 128
rect 52 240 88 248
rect 52 128 60 240
rect 80 128 88 240
rect 52 120 88 128
rect 112 240 148 248
rect 112 128 120 240
rect 140 128 148 240
rect 176 240 212 248
rect 176 152 184 240
rect 204 152 212 240
rect 176 144 212 152
rect 236 240 272 248
rect 236 152 244 240
rect 264 152 272 240
rect 236 144 272 152
rect 300 240 336 248
rect 300 152 308 240
rect 328 152 336 240
rect 300 144 336 152
rect 360 240 396 248
rect 360 152 368 240
rect 388 152 396 240
rect 360 144 396 152
rect 112 120 148 128
rect 204 116 244 124
rect -44 92 -4 100
rect -44 68 -36 92
rect -12 68 -4 92
rect -44 60 -4 68
rect 80 92 120 100
rect 80 68 88 92
rect 112 68 120 92
rect 204 92 212 116
rect 236 92 244 116
rect 204 84 244 92
rect 328 116 368 124
rect 328 92 336 116
rect 360 92 368 116
rect 328 84 368 92
rect 80 60 120 68
rect 176 56 212 64
rect -128 28 -92 36
rect -24 28 12 36
rect -128 8 -120 28
rect -100 8 -16 28
rect 4 8 12 28
rect -128 0 -92 8
rect -24 0 12 8
rect 80 28 120 36
rect 80 4 88 28
rect 112 4 120 28
rect 176 20 184 56
rect 204 20 212 56
rect 176 12 212 20
rect 236 56 272 64
rect 236 20 244 56
rect 264 20 272 56
rect 236 12 272 20
rect 300 56 336 64
rect 300 20 308 56
rect 328 20 336 56
rect 300 12 336 20
rect 360 56 396 64
rect 360 20 368 56
rect 388 20 396 56
rect 360 12 396 20
rect 80 -4 120 4
rect -72 -32 -36 -24
rect -72 -196 -64 -32
rect -44 -196 -36 -32
rect -72 -204 -36 -196
rect -12 -32 24 -24
rect -12 -196 -4 -32
rect 16 -196 24 -32
rect -12 -204 24 -196
rect 52 -32 88 -24
rect 52 -196 60 -32
rect 80 -196 88 -32
rect 52 -204 88 -196
rect 112 -32 148 -24
rect 112 -196 120 -32
rect 140 -196 148 -32
rect 204 -60 244 -52
rect 328 -60 368 -52
rect 204 -84 212 -60
rect 236 -80 336 -60
rect 236 -84 244 -80
rect 204 -92 244 -84
rect 328 -84 336 -80
rect 360 -84 368 -60
rect 328 -92 368 -84
rect 112 -204 148 -196
rect 176 -120 212 -112
rect 176 -196 184 -120
rect 204 -196 212 -120
rect 176 -204 212 -196
rect 236 -120 272 -112
rect 236 -196 244 -120
rect 264 -196 272 -120
rect 236 -204 272 -196
rect 300 -120 336 -112
rect 300 -196 308 -120
rect 328 -196 336 -120
rect 300 -204 336 -196
rect 360 -120 396 -112
rect 360 -196 368 -120
rect 388 -196 396 -120
rect 360 -204 396 -196
rect -44 -232 -4 -224
rect -44 -256 -36 -232
rect -12 -256 -4 -232
rect -44 -264 -4 -256
rect -88 -320 -28 -300
rect -88 -340 -68 -320
rect -48 -340 -28 -320
rect -88 -360 -28 -340
<< viali >>
rect 36 284 56 304
rect 460 284 480 304
rect -64 128 -44 240
rect -4 128 16 240
rect 60 128 80 240
rect 120 128 140 240
rect 184 152 204 240
rect 244 152 264 240
rect 308 152 328 240
rect 368 152 388 240
rect -36 68 -12 92
rect 88 68 112 92
rect 212 92 236 116
rect 336 92 360 116
rect -120 8 -100 28
rect -16 8 4 28
rect 88 4 112 28
rect 184 20 204 56
rect 244 20 264 56
rect 308 20 328 56
rect 368 20 388 56
rect -64 -196 -44 -32
rect -4 -196 16 -32
rect 60 -196 80 -32
rect 120 -196 140 -32
rect 212 -84 236 -60
rect 336 -84 360 -60
rect 184 -196 204 -120
rect 244 -196 264 -120
rect 308 -196 328 -120
rect 368 -196 388 -120
rect -36 -256 -12 -232
rect 368 -296 388 -276
rect -68 -340 -48 -320
<< metal1 >>
rect 4 312 88 324
rect -140 304 488 312
rect -140 284 36 304
rect 56 284 460 304
rect 480 284 488 304
rect -140 276 488 284
rect -140 268 452 276
rect -72 240 -36 248
rect -72 128 -64 240
rect -44 128 -36 240
rect -72 120 -36 128
rect -12 240 24 268
rect -12 128 -4 240
rect 16 128 24 240
rect -12 120 24 128
rect 52 240 88 268
rect 52 128 60 240
rect 80 128 88 240
rect 52 120 88 128
rect 112 240 148 248
rect 112 128 120 240
rect 140 128 148 240
rect 176 240 212 268
rect 176 152 184 240
rect 204 152 212 240
rect 176 144 212 152
rect 236 240 272 248
rect 236 152 244 240
rect 264 156 272 240
rect 300 240 336 268
rect 264 152 276 156
rect 236 144 276 152
rect 300 152 308 240
rect 328 152 336 240
rect 300 144 336 152
rect 360 240 396 248
rect 360 152 368 240
rect 388 156 396 240
rect 388 152 400 156
rect 360 144 400 152
rect 112 120 152 128
rect -72 100 -44 120
rect 136 112 152 120
rect 204 116 244 124
rect 204 112 212 116
rect -72 92 -4 100
rect -72 68 -36 92
rect -12 88 -4 92
rect 80 92 120 100
rect 80 88 88 92
rect -12 72 88 88
rect -12 68 -4 72
rect -72 60 -4 68
rect 80 68 88 72
rect 112 68 120 92
rect 80 60 120 68
rect 136 96 212 112
rect -128 28 -92 36
rect -128 8 -120 28
rect -100 8 -92 28
rect -128 0 -92 8
rect -72 -24 -44 60
rect -24 28 12 36
rect -24 8 -16 28
rect 4 24 12 28
rect 80 28 120 36
rect 80 24 88 28
rect 4 8 88 24
rect -24 0 12 8
rect 80 4 88 8
rect 112 4 120 28
rect 80 -4 120 4
rect 136 -24 152 96
rect 204 92 212 96
rect 236 92 244 116
rect 204 84 244 92
rect 260 112 276 144
rect 328 116 368 124
rect 328 112 336 116
rect 260 96 336 112
rect 260 64 276 96
rect 328 92 336 96
rect 360 92 368 116
rect 328 84 368 92
rect 384 112 400 144
rect 384 96 524 112
rect 384 64 400 96
rect 176 56 212 64
rect 176 20 184 56
rect 204 20 212 56
rect 176 12 212 20
rect 236 56 276 64
rect 236 20 244 56
rect 264 52 276 56
rect 300 56 336 64
rect 264 20 272 52
rect 236 12 272 20
rect 300 20 308 56
rect 328 20 336 56
rect 300 12 336 20
rect 360 56 400 64
rect 360 20 368 56
rect 388 52 400 56
rect 388 20 396 52
rect 360 12 396 20
rect 176 -8 192 12
rect 300 -8 316 12
rect 176 -24 316 -8
rect -72 -32 -36 -24
rect -72 -196 -64 -32
rect -44 -196 -36 -32
rect -72 -204 -36 -196
rect -12 -32 24 -24
rect -12 -196 -4 -32
rect 16 -184 24 -32
rect 52 -32 88 -24
rect 52 -184 60 -32
rect 16 -196 60 -184
rect 80 -196 88 -32
rect -12 -204 88 -196
rect 112 -32 152 -24
rect 112 -196 120 -32
rect 140 -36 152 -32
rect 140 -196 148 -36
rect 204 -60 244 -52
rect 204 -84 212 -60
rect 236 -84 244 -60
rect 204 -92 244 -84
rect 272 -112 300 -24
rect 328 -60 396 -52
rect 328 -84 336 -60
rect 360 -84 396 -60
rect 328 -92 396 -84
rect 368 -112 396 -92
rect 112 -204 148 -196
rect 176 -120 212 -112
rect 176 -196 184 -120
rect 204 -196 212 -120
rect 176 -204 212 -196
rect 236 -120 336 -112
rect 236 -196 244 -120
rect 264 -128 308 -120
rect 264 -184 272 -128
rect 300 -184 308 -128
rect 264 -196 308 -184
rect 328 -196 336 -120
rect 236 -204 336 -196
rect 360 -120 396 -112
rect 360 -196 368 -120
rect 388 -196 396 -120
rect 52 -224 68 -204
rect 176 -224 200 -204
rect -44 -232 -4 -224
rect -44 -236 -36 -232
rect -100 -252 -36 -236
rect -44 -256 -36 -252
rect -12 -256 -4 -232
rect 52 -240 200 -224
rect -44 -264 -4 -256
rect -88 -320 -28 -300
rect 272 -320 300 -204
rect 360 -276 396 -196
rect 360 -296 368 -276
rect 388 -296 396 -276
rect 360 -304 396 -296
rect -140 -340 -68 -320
rect -48 -340 452 -320
rect -140 -360 452 -340
<< labels >>
rlabel metal1 268 100 276 104 1 vinv
port 6 n
rlabel metal1 392 100 400 104 1 vout
port 1 n
rlabel metal1 -116 4 -108 8 1 vin2
port 4 n
rlabel metal1 -80 -248 -72 -244 1 vin1
port 3 n
rlabel metal1 32 72 40 76 1 vg34
rlabel metal1 144 32 152 36 1 vamp
port 7 n
rlabel metal1 116 -236 124 -232 1 vs12
rlabel metal1 380 -224 388 -220 1 Vtail
rlabel metal1 104 -348 112 -340 1 gnd
port 2 n
rlabel metal1 -88 292 -80 296 1 vdd
port 5 n
<< end >>
