magic
tech sky130A
timestamp 1762235650
<< nwell >>
rect -100 -20 100 160
<< pmos >>
rect -10 0 10 140
<< pdiff >>
rect -80 130 -10 140
rect -80 10 -70 130
rect -50 10 -10 130
rect -80 0 -10 10
rect 10 130 80 140
rect 10 10 50 130
rect 70 10 80 130
rect 10 0 80 10
<< pdiffc >>
rect -70 10 -50 130
rect 50 10 70 130
<< poly >>
rect -10 140 10 160
rect -10 -20 10 0
<< locali >>
rect -80 130 -40 140
rect -80 10 -70 130
rect -50 10 -40 130
rect -80 0 -40 10
rect 40 130 80 140
rect 40 10 50 130
rect 70 10 80 130
rect 40 0 80 10
<< end >>
