magic
tech sky130A
timestamp 1764654977
<< nwell >>
rect 40 230 150 310
rect -100 30 680 230
rect 270 -20 680 30
<< nmos >>
rect -20 -220 20 -100
rect 170 -220 210 -100
rect 370 -130 410 -80
rect 560 -130 600 -80
rect 100 -420 140 -350
rect 290 -420 330 -350
<< pmos >>
rect -20 50 20 210
rect 170 50 210 210
rect 370 0 410 210
rect 560 0 600 210
<< ndiff >>
rect 310 -90 370 -80
rect -80 -110 -20 -100
rect -80 -210 -70 -110
rect -50 -210 -20 -110
rect -80 -220 -20 -210
rect 20 -110 80 -100
rect 20 -210 50 -110
rect 70 -210 80 -110
rect 20 -220 80 -210
rect 110 -110 170 -100
rect 110 -210 120 -110
rect 140 -210 170 -110
rect 110 -220 170 -210
rect 210 -110 270 -100
rect 210 -210 240 -110
rect 260 -210 270 -110
rect 310 -120 320 -90
rect 340 -120 370 -90
rect 310 -130 370 -120
rect 410 -90 470 -80
rect 410 -120 440 -90
rect 460 -120 470 -90
rect 410 -130 470 -120
rect 500 -90 560 -80
rect 500 -120 510 -90
rect 530 -120 560 -90
rect 500 -130 560 -120
rect 600 -90 660 -80
rect 600 -120 630 -90
rect 650 -120 660 -90
rect 600 -130 660 -120
rect 210 -220 270 -210
rect 40 -360 100 -350
rect 40 -410 50 -360
rect 70 -410 100 -360
rect 40 -420 100 -410
rect 140 -360 200 -350
rect 140 -410 170 -360
rect 190 -410 200 -360
rect 140 -420 200 -410
rect 230 -360 290 -350
rect 230 -410 240 -360
rect 260 -410 290 -360
rect 230 -420 290 -410
rect 330 -360 390 -350
rect 330 -410 360 -360
rect 380 -410 390 -360
rect 330 -420 390 -410
<< pdiff >>
rect -80 200 -20 210
rect -80 60 -70 200
rect -50 60 -20 200
rect -80 50 -20 60
rect 20 200 80 210
rect 20 60 50 200
rect 70 60 80 200
rect 20 50 80 60
rect 110 200 170 210
rect 110 60 120 200
rect 140 60 170 200
rect 110 50 170 60
rect 210 200 270 210
rect 210 60 240 200
rect 260 60 270 200
rect 210 50 270 60
rect 310 200 370 210
rect 310 10 320 200
rect 340 10 370 200
rect 310 0 370 10
rect 410 200 470 210
rect 410 10 440 200
rect 460 10 470 200
rect 410 0 470 10
rect 500 200 560 210
rect 500 10 510 200
rect 530 10 560 200
rect 500 0 560 10
rect 600 200 660 210
rect 600 10 630 200
rect 650 10 660 200
rect 600 0 660 10
<< ndiffc >>
rect -70 -210 -50 -110
rect 50 -210 70 -110
rect 120 -210 140 -110
rect 240 -210 260 -110
rect 320 -120 340 -90
rect 440 -120 460 -90
rect 510 -120 530 -90
rect 630 -120 650 -90
rect 50 -410 70 -360
rect 170 -410 190 -360
rect 240 -410 260 -360
rect 360 -410 380 -360
<< pdiffc >>
rect -70 60 -50 200
rect 50 60 70 200
rect 120 60 140 200
rect 240 60 260 200
rect 320 10 340 200
rect 440 10 460 200
rect 510 10 530 200
rect 630 10 650 200
<< psubdiff >>
rect -100 -380 -40 -360
rect -100 -400 -80 -380
rect -60 -400 -40 -380
rect -100 -420 -40 -400
<< nsubdiff >>
rect 75 275 115 290
rect 75 255 85 275
rect 105 255 115 275
rect 75 240 115 255
<< psubdiffcont >>
rect -80 -400 -60 -380
<< nsubdiffcont >>
rect 85 255 105 275
<< poly >>
rect -20 210 20 240
rect 170 210 210 240
rect 370 210 410 240
rect 560 210 600 240
rect -20 20 20 50
rect -20 0 -10 20
rect 10 0 20 20
rect -20 -10 20 0
rect 170 20 210 50
rect 170 0 180 20
rect 200 0 210 20
rect 170 -10 210 0
rect 370 -30 410 0
rect 170 -50 210 -40
rect 170 -70 180 -50
rect 200 -70 210 -50
rect -20 -100 20 -80
rect 170 -100 210 -70
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -80 410 -50
rect 560 -30 600 0
rect 560 -50 570 -30
rect 590 -50 600 -30
rect 560 -80 600 -50
rect 370 -150 410 -130
rect 560 -150 600 -130
rect -20 -249 20 -220
rect 170 -240 210 -220
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 100 -300 140 -290
rect 100 -320 110 -300
rect 130 -320 140 -300
rect 100 -350 140 -320
rect 290 -300 330 -290
rect 290 -320 300 -300
rect 320 -320 330 -300
rect 290 -350 330 -320
rect 100 -440 140 -420
rect 290 -440 330 -420
<< polycont >>
rect -10 0 10 20
rect 180 0 200 20
rect 180 -70 200 -50
rect 380 -50 400 -30
rect 570 -50 590 -30
rect -11 -269 10 -249
rect 110 -320 130 -300
rect 300 -320 320 -300
<< xpolycontact >>
rect 720 -290 760 30
rect 440 -330 660 -290
<< xpolyres >>
rect 660 -330 760 -290
<< locali >>
rect 720 300 760 310
rect 75 275 115 285
rect 75 255 85 275
rect 105 255 115 275
rect 75 245 115 255
rect 720 280 730 300
rect 750 280 760 300
rect -80 200 -40 210
rect -80 60 -70 200
rect -50 60 -40 200
rect -80 50 -40 60
rect 40 200 80 210
rect 40 60 50 200
rect 70 60 80 200
rect 40 50 80 60
rect 110 200 150 210
rect 110 60 120 200
rect 140 60 150 200
rect 110 50 150 60
rect 230 200 270 210
rect 230 60 240 200
rect 260 60 270 200
rect 230 50 270 60
rect 310 200 350 210
rect -20 20 20 30
rect -20 0 -10 20
rect 10 0 20 20
rect -20 -10 20 0
rect 170 20 210 30
rect 170 0 180 20
rect 200 0 210 20
rect 310 10 320 200
rect 340 10 350 200
rect 310 0 350 10
rect 430 200 470 210
rect 430 10 440 200
rect 460 10 470 200
rect 430 0 470 10
rect 500 200 540 210
rect 500 10 510 200
rect 530 10 540 200
rect 500 0 540 10
rect 620 200 660 210
rect 620 10 630 200
rect 650 10 660 200
rect 720 180 760 280
rect 720 160 730 180
rect 750 160 760 180
rect 720 150 760 160
rect 620 0 660 10
rect 170 -10 210 0
rect 370 -30 410 -20
rect -140 -50 20 -40
rect -140 -70 -130 -50
rect -110 -70 -10 -50
rect 10 -70 20 -50
rect -140 -80 20 -70
rect 170 -50 210 -40
rect 170 -70 180 -50
rect 200 -70 210 -50
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -60 410 -50
rect 560 -30 600 -20
rect 560 -50 570 -30
rect 590 -50 600 -30
rect 560 -60 600 -50
rect 170 -80 210 -70
rect 310 -90 350 -80
rect -80 -110 -40 -100
rect -80 -210 -70 -110
rect -50 -210 -40 -110
rect -80 -220 -40 -210
rect 40 -110 80 -100
rect 40 -210 50 -110
rect 70 -210 80 -110
rect 40 -220 80 -210
rect 110 -110 150 -100
rect 110 -210 120 -110
rect 140 -210 150 -110
rect 110 -220 150 -210
rect 230 -110 270 -100
rect 230 -210 240 -110
rect 260 -210 270 -110
rect 310 -120 320 -90
rect 340 -120 350 -90
rect 310 -130 350 -120
rect 430 -90 470 -80
rect 430 -120 440 -90
rect 460 -120 470 -90
rect 430 -130 470 -120
rect 500 -90 540 -80
rect 500 -120 510 -90
rect 530 -120 540 -90
rect 500 -130 540 -120
rect 620 -90 660 -80
rect 620 -120 630 -90
rect 650 -120 660 -90
rect 620 -130 660 -120
rect 230 -220 270 -210
rect -20 -249 20 -240
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 100 -300 140 -290
rect 100 -320 110 -300
rect 130 -320 140 -300
rect 100 -330 140 -320
rect 290 -300 330 -290
rect 290 -320 300 -300
rect 320 -320 330 -300
rect 290 -330 330 -320
rect 40 -360 80 -350
rect -100 -380 -40 -360
rect -100 -400 -80 -380
rect -60 -400 -40 -380
rect -100 -420 -40 -400
rect 40 -410 50 -360
rect 70 -410 80 -360
rect 40 -420 80 -410
rect 160 -360 200 -350
rect 160 -410 170 -360
rect 190 -410 200 -360
rect 160 -420 200 -410
rect 230 -360 270 -350
rect 230 -410 240 -360
rect 260 -410 270 -360
rect 230 -420 270 -410
rect 350 -360 390 -350
rect 350 -410 360 -360
rect 380 -410 390 -360
rect 350 -420 390 -410
<< viali >>
rect 85 255 105 275
rect 730 280 750 300
rect -70 60 -50 200
rect 50 60 70 200
rect 120 60 140 200
rect 240 60 260 200
rect -10 0 10 20
rect 180 0 200 20
rect 320 10 340 200
rect 440 10 460 200
rect 510 10 530 200
rect 630 10 650 200
rect 730 160 750 180
rect 730 0 750 20
rect -130 -70 -110 -50
rect -10 -70 10 -50
rect 180 -70 200 -50
rect 380 -50 400 -30
rect 570 -50 590 -30
rect -70 -210 -50 -110
rect 50 -210 70 -110
rect 120 -210 140 -110
rect 240 -210 260 -110
rect 320 -120 340 -90
rect 440 -120 460 -90
rect 510 -120 530 -90
rect 630 -120 650 -90
rect -11 -269 10 -249
rect 110 -320 130 -300
rect 300 -320 320 -300
rect 450 -320 470 -300
rect -80 -400 -60 -380
rect 50 -410 70 -360
rect 170 -410 190 -360
rect 240 -410 260 -360
rect 360 -410 380 -360
<< metal1 >>
rect -140 300 760 310
rect -140 280 730 300
rect 750 280 760 300
rect -140 275 760 280
rect -140 270 85 275
rect 40 255 85 270
rect 105 270 760 275
rect 105 255 150 270
rect 40 230 150 255
rect -80 200 -40 210
rect -80 60 -70 200
rect -50 60 -40 200
rect -80 30 -40 60
rect 40 200 80 230
rect 40 60 50 200
rect 70 60 80 200
rect 40 50 80 60
rect 110 200 150 230
rect 110 60 120 200
rect 140 60 150 200
rect 110 50 150 60
rect 230 200 270 210
rect 230 60 240 200
rect 260 60 270 200
rect -80 20 210 30
rect -80 0 -10 20
rect 10 0 180 20
rect 200 0 210 20
rect -80 -10 210 0
rect -140 -50 -100 -40
rect -140 -70 -130 -50
rect -110 -70 -100 -50
rect -140 -80 -100 -70
rect -80 -110 -40 -10
rect 230 -20 270 60
rect 310 200 350 270
rect 310 10 320 200
rect 340 10 350 200
rect 310 0 350 10
rect 430 200 470 210
rect 430 10 440 200
rect 460 10 470 200
rect 230 -30 410 -20
rect -20 -50 210 -40
rect -20 -70 -10 -50
rect 10 -70 180 -50
rect 200 -70 210 -50
rect -20 -80 210 -70
rect 230 -50 380 -30
rect 400 -50 410 -30
rect 230 -60 410 -50
rect 430 -21 470 10
rect 500 200 540 270
rect 500 10 510 200
rect 530 10 540 200
rect 500 0 540 10
rect 620 210 830 250
rect 620 200 660 210
rect 620 10 630 200
rect 650 10 660 200
rect 500 -21 600 -20
rect 430 -30 600 -21
rect 430 -50 570 -30
rect 590 -50 600 -30
rect 430 -60 600 -50
rect -80 -210 -70 -110
rect -50 -210 -40 -110
rect -80 -220 -40 -210
rect 40 -110 80 -100
rect 40 -210 50 -110
rect 70 -210 80 -110
rect 110 -110 150 -100
rect 110 -210 120 -110
rect 140 -210 150 -110
rect -140 -249 20 -240
rect -140 -269 -11 -249
rect 10 -269 20 -249
rect -140 -280 20 -269
rect 40 -260 150 -210
rect 230 -110 270 -60
rect 230 -210 240 -110
rect 260 -210 270 -110
rect 230 -220 270 -210
rect 310 -90 350 -80
rect 310 -120 320 -90
rect 340 -120 350 -90
rect 310 -230 350 -120
rect 430 -90 470 -60
rect 430 -120 440 -90
rect 460 -120 470 -90
rect 430 -130 470 -120
rect 500 -90 540 -80
rect 500 -120 510 -90
rect 530 -120 540 -90
rect 500 -230 540 -120
rect 620 -90 660 10
rect 720 180 760 190
rect 720 160 730 180
rect 750 160 760 180
rect 720 20 760 160
rect 720 0 730 20
rect 750 0 760 20
rect 720 -10 760 0
rect 620 -120 630 -90
rect 650 -120 660 -90
rect 620 -130 660 -120
rect 40 -360 80 -260
rect 310 -270 540 -230
rect 100 -300 480 -290
rect 100 -320 110 -300
rect 130 -320 300 -300
rect 320 -320 450 -300
rect 470 -320 480 -300
rect 100 -330 480 -320
rect -100 -380 -40 -360
rect -100 -400 -80 -380
rect -60 -400 -40 -380
rect -100 -460 -40 -400
rect 40 -410 50 -360
rect 70 -410 80 -360
rect 40 -420 80 -410
rect 160 -360 200 -350
rect 160 -410 170 -360
rect 190 -410 200 -360
rect 160 -460 200 -410
rect 230 -360 270 -350
rect 230 -410 240 -360
rect 260 -410 270 -360
rect 230 -460 270 -410
rect 350 -360 390 -330
rect 350 -410 360 -360
rect 380 -410 390 -360
rect 350 -420 390 -410
rect 500 -460 540 -270
rect -140 -500 540 -460
<< labels >>
rlabel metal1 -65 305 -64 306 1 Vdd
rlabel metal1 322 -45 334 -35 1 vinv
rlabel metal1 460 -50 480 -30 1 vinv2
rlabel metal1 90 -230 90 -230 1 VS12
rlabel metal1 -61 -261 -57 -255 1 vin1
rlabel metal1 55 10 55 10 1 VG34
rlabel viali -120 -60 -120 -60 1 vin2
rlabel metal1 170 -490 200 -480 1 Gnd
rlabel metal1 800 220 820 240 1 vout
<< end >>
