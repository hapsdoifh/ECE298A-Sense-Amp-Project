magic
tech sky130A
timestamp 1764712608
<< nwell >>
rect 40 230 150 310
rect -100 130 680 230
rect 270 90 680 130
<< nmos >>
rect -20 -190 20 -10
rect 170 -190 210 -10
rect 370 -20 410 30
rect 560 -20 600 30
rect 370 -260 410 -170
rect 560 -260 600 -170
<< pmos >>
rect -20 150 20 210
rect 170 150 210 210
rect 370 110 410 210
rect 560 110 600 210
<< ndiff >>
rect 310 20 370 30
rect 310 -10 320 20
rect 340 -10 370 20
rect -80 -20 -20 -10
rect -80 -180 -70 -20
rect -50 -180 -20 -20
rect -80 -190 -20 -180
rect 20 -20 80 -10
rect 20 -180 50 -20
rect 70 -180 80 -20
rect 20 -190 80 -180
rect 110 -20 170 -10
rect 110 -180 120 -20
rect 140 -180 170 -20
rect 110 -190 170 -180
rect 210 -20 270 -10
rect 310 -20 370 -10
rect 410 20 470 30
rect 410 -10 440 20
rect 460 -10 470 20
rect 410 -20 470 -10
rect 500 20 560 30
rect 500 -10 510 20
rect 530 -10 560 20
rect 500 -20 560 -10
rect 600 20 660 30
rect 600 -10 630 20
rect 650 -10 660 20
rect 600 -20 660 -10
rect 210 -180 240 -20
rect 260 -180 270 -20
rect 210 -190 270 -180
rect 310 -180 370 -170
rect 310 -250 320 -180
rect 340 -250 370 -180
rect 310 -260 370 -250
rect 410 -180 470 -170
rect 410 -250 440 -180
rect 460 -250 470 -180
rect 410 -260 470 -250
rect 500 -180 560 -170
rect 500 -250 510 -180
rect 530 -250 560 -180
rect 500 -260 560 -250
rect 600 -180 660 -170
rect 600 -250 630 -180
rect 650 -250 660 -180
rect 600 -260 660 -250
<< pdiff >>
rect -80 200 -20 210
rect -80 160 -70 200
rect -50 160 -20 200
rect -80 150 -20 160
rect 20 200 80 210
rect 20 160 50 200
rect 70 160 80 200
rect 20 150 80 160
rect 110 200 170 210
rect 110 160 120 200
rect 140 160 170 200
rect 110 150 170 160
rect 210 200 270 210
rect 210 160 240 200
rect 260 160 270 200
rect 210 150 270 160
rect 310 200 370 210
rect 310 120 320 200
rect 340 120 370 200
rect 310 110 370 120
rect 410 200 470 210
rect 410 120 440 200
rect 460 120 470 200
rect 410 110 470 120
rect 500 200 560 210
rect 500 120 510 200
rect 530 120 560 200
rect 500 110 560 120
rect 600 200 660 210
rect 600 120 630 200
rect 650 120 660 200
rect 600 110 660 120
<< ndiffc >>
rect 320 -10 340 20
rect -70 -180 -50 -20
rect 50 -180 70 -20
rect 120 -180 140 -20
rect 440 -10 460 20
rect 510 -10 530 20
rect 630 -10 650 20
rect 240 -180 260 -20
rect 320 -250 340 -180
rect 440 -250 460 -180
rect 510 -250 530 -180
rect 630 -250 650 -180
<< pdiffc >>
rect -70 160 -50 200
rect 50 160 70 200
rect 120 160 140 200
rect 240 160 260 200
rect 320 120 340 200
rect 440 120 460 200
rect 510 120 530 200
rect 630 120 650 200
<< psubdiff >>
rect 40 -300 100 -280
rect 40 -320 60 -300
rect 80 -320 100 -300
rect 40 -340 100 -320
<< nsubdiff >>
rect 75 275 115 290
rect 75 255 85 275
rect 105 255 115 275
rect 75 240 115 255
<< psubdiffcont >>
rect 60 -320 80 -300
<< nsubdiffcont >>
rect 85 255 105 275
<< poly >>
rect -20 210 20 240
rect 170 210 210 240
rect 370 210 410 240
rect 560 210 600 240
rect -20 120 20 150
rect -20 100 -10 120
rect 10 100 20 120
rect -20 90 20 100
rect 170 120 210 150
rect 170 100 180 120
rect 200 100 210 120
rect 170 90 210 100
rect 370 80 410 110
rect 370 60 380 80
rect 400 60 410 80
rect 170 40 210 50
rect 170 20 180 40
rect 200 20 210 40
rect 370 30 410 60
rect 560 80 600 110
rect 560 60 570 80
rect 590 60 600 80
rect 560 30 600 60
rect -20 -10 20 10
rect 170 -10 210 20
rect 370 -40 410 -20
rect 560 -40 600 -20
rect 370 -120 410 -110
rect 370 -140 380 -120
rect 400 -140 410 -120
rect 370 -170 410 -140
rect 560 -120 600 -110
rect 560 -140 570 -120
rect 590 -140 600 -120
rect 560 -170 600 -140
rect -20 -219 20 -190
rect 170 -210 210 -190
rect -20 -239 -11 -219
rect 10 -239 20 -219
rect -20 -250 20 -239
rect 370 -280 410 -260
rect 560 -280 600 -260
<< polycont >>
rect -10 100 10 120
rect 180 100 200 120
rect 380 60 400 80
rect 180 20 200 40
rect 570 60 590 80
rect 380 -140 400 -120
rect 570 -140 590 -120
rect -11 -239 10 -219
<< xpolycontact >>
rect 720 90 760 310
rect 720 -210 760 10
<< xpolyres >>
rect 720 10 760 90
<< locali >>
rect 75 275 115 285
rect 75 255 85 275
rect 105 255 115 275
rect 75 245 115 255
rect -80 200 -40 210
rect -80 160 -70 200
rect -50 160 -40 200
rect -80 150 -40 160
rect 40 200 80 210
rect 40 160 50 200
rect 70 160 80 200
rect 40 150 80 160
rect 110 200 150 210
rect 110 160 120 200
rect 140 160 150 200
rect 110 150 150 160
rect 230 200 270 210
rect 230 160 240 200
rect 260 160 270 200
rect 230 150 270 160
rect 310 200 350 210
rect -20 120 20 130
rect -20 100 -10 120
rect 10 100 20 120
rect -20 90 20 100
rect 170 120 210 130
rect 170 100 180 120
rect 200 100 210 120
rect 310 120 320 200
rect 340 120 350 200
rect 310 110 350 120
rect 430 200 470 210
rect 430 120 440 200
rect 460 120 470 200
rect 430 110 470 120
rect 500 200 540 210
rect 500 120 510 200
rect 530 120 540 200
rect 500 110 540 120
rect 620 200 660 210
rect 620 120 630 200
rect 650 120 660 200
rect 620 110 660 120
rect 170 90 210 100
rect 370 80 410 90
rect 370 60 380 80
rect 400 60 410 80
rect 370 50 410 60
rect 560 80 600 90
rect 560 60 570 80
rect 590 60 600 80
rect 560 50 600 60
rect -140 40 20 50
rect -140 20 -130 40
rect -110 20 -10 40
rect 10 20 20 40
rect -140 10 20 20
rect 170 40 210 50
rect 170 20 180 40
rect 200 20 210 40
rect 170 10 210 20
rect 310 20 350 30
rect 310 -10 320 20
rect 340 -10 350 20
rect -80 -20 -40 -10
rect -80 -180 -70 -20
rect -50 -180 -40 -20
rect -80 -190 -40 -180
rect 40 -20 80 -10
rect 40 -180 50 -20
rect 70 -180 80 -20
rect 40 -190 80 -180
rect 110 -20 150 -10
rect 110 -180 120 -20
rect 140 -180 150 -20
rect 110 -190 150 -180
rect 230 -20 270 -10
rect 310 -20 350 -10
rect 430 20 470 30
rect 430 -10 440 20
rect 460 -10 470 20
rect 430 -20 470 -10
rect 500 20 540 30
rect 500 -10 510 20
rect 530 -10 540 20
rect 500 -20 540 -10
rect 620 20 660 30
rect 620 -10 630 20
rect 650 -10 660 20
rect 620 -20 660 -10
rect 230 -180 240 -20
rect 260 -180 270 -20
rect 500 -60 540 -50
rect 500 -80 510 -60
rect 530 -80 540 -60
rect 370 -120 410 -110
rect 370 -140 380 -120
rect 400 -140 410 -120
rect 370 -150 410 -140
rect 230 -190 270 -180
rect 310 -180 350 -170
rect -20 -219 20 -210
rect -20 -239 -11 -219
rect 10 -239 20 -219
rect -20 -250 20 -239
rect 310 -250 320 -180
rect 340 -250 350 -180
rect 310 -260 350 -250
rect 430 -180 470 -170
rect 430 -250 440 -180
rect 460 -250 470 -180
rect 430 -260 470 -250
rect 500 -180 540 -80
rect 560 -120 600 -110
rect 560 -140 570 -120
rect 590 -140 600 -120
rect 560 -150 600 -140
rect 500 -250 510 -180
rect 530 -250 540 -180
rect 500 -260 540 -250
rect 620 -180 660 -170
rect 620 -250 630 -180
rect 650 -250 660 -180
rect 620 -260 660 -250
rect 40 -300 100 -280
rect 40 -320 60 -300
rect 80 -320 100 -300
rect 40 -340 100 -320
<< viali >>
rect 85 255 105 275
rect 730 280 750 300
rect -70 160 -50 200
rect 50 160 70 200
rect 120 160 140 200
rect 240 160 260 200
rect -10 100 10 120
rect 180 100 200 120
rect 320 120 340 200
rect 440 120 460 200
rect 510 120 530 200
rect 630 120 650 200
rect 380 60 400 80
rect 570 60 590 80
rect -130 20 -110 40
rect -10 20 10 40
rect 180 20 200 40
rect 320 -10 340 20
rect -70 -180 -50 -20
rect 50 -180 70 -20
rect 120 -180 140 -20
rect 440 -10 460 20
rect 510 -10 530 20
rect 630 -10 650 20
rect 240 -180 260 -20
rect 510 -80 530 -60
rect 380 -140 400 -120
rect -11 -239 10 -219
rect 320 -250 340 -180
rect 440 -250 460 -180
rect 570 -140 590 -120
rect 510 -250 530 -180
rect 630 -250 650 -180
rect 730 -200 750 -180
rect 60 -320 80 -300
<< metal1 >>
rect -140 300 760 310
rect -140 280 730 300
rect 750 280 760 300
rect -140 275 760 280
rect -140 270 85 275
rect 40 255 85 270
rect 105 270 760 275
rect 105 255 150 270
rect 40 230 150 255
rect -80 200 -40 210
rect -80 160 -70 200
rect -50 160 -40 200
rect -80 130 -40 160
rect 40 200 80 230
rect 40 160 50 200
rect 70 160 80 200
rect 40 150 80 160
rect 110 200 150 230
rect 110 160 120 200
rect 140 160 150 200
rect 110 150 150 160
rect 230 200 270 210
rect 230 160 240 200
rect 260 160 270 200
rect -80 120 210 130
rect -80 100 -10 120
rect 10 100 180 120
rect 200 100 210 120
rect -80 90 210 100
rect 230 90 270 160
rect 310 200 350 270
rect 310 120 320 200
rect 340 120 350 200
rect 310 110 350 120
rect 430 200 470 210
rect 430 120 440 200
rect 460 120 470 200
rect -140 40 -100 50
rect -140 20 -130 40
rect -110 20 -100 40
rect -140 10 -100 20
rect -80 -20 -40 90
rect 230 80 410 90
rect 230 60 380 80
rect 400 60 410 80
rect 230 50 410 60
rect 430 89 470 120
rect 500 200 540 270
rect 500 120 510 200
rect 530 120 540 200
rect 500 110 540 120
rect 620 210 830 250
rect 620 200 660 210
rect 620 120 630 200
rect 650 120 660 200
rect 500 89 600 90
rect 430 80 600 89
rect 430 60 570 80
rect 590 60 600 80
rect 430 50 600 60
rect -20 40 210 50
rect -20 20 -10 40
rect 10 20 180 40
rect 200 20 210 40
rect -20 10 210 20
rect -80 -180 -70 -20
rect -50 -180 -40 -20
rect -80 -190 -40 -180
rect 40 -20 80 -10
rect 40 -180 50 -20
rect 70 -150 80 -20
rect 110 -20 150 -10
rect 110 -150 120 -20
rect 70 -180 120 -150
rect 140 -180 150 -20
rect 40 -190 150 -180
rect 230 -20 270 50
rect 230 -180 240 -20
rect 260 -180 270 -20
rect 310 20 350 30
rect 310 -10 320 20
rect 340 -10 350 20
rect 310 -50 350 -10
rect 430 20 470 50
rect 430 -10 440 20
rect 460 -10 470 20
rect 430 -20 470 -10
rect 500 20 540 30
rect 500 -10 510 20
rect 530 -10 540 20
rect 500 -50 540 -10
rect 620 20 660 120
rect 620 -10 630 20
rect 650 -10 660 20
rect 620 -20 660 -10
rect 310 -60 540 -50
rect 310 -80 510 -60
rect 530 -80 540 -60
rect 310 -90 540 -80
rect 370 -120 660 -110
rect 370 -140 380 -120
rect 400 -140 570 -120
rect 590 -140 660 -120
rect 370 -150 660 -140
rect 620 -170 660 -150
rect 230 -190 270 -180
rect 310 -180 350 -170
rect -140 -219 20 -210
rect -140 -239 -11 -219
rect 10 -239 20 -219
rect -140 -250 20 -239
rect 110 -220 150 -190
rect 310 -220 320 -180
rect 110 -250 320 -220
rect 340 -250 350 -180
rect 110 -260 350 -250
rect 430 -180 470 -170
rect 430 -250 440 -180
rect 460 -250 470 -180
rect 40 -300 100 -280
rect 430 -300 470 -250
rect 500 -180 540 -170
rect 500 -250 510 -180
rect 530 -250 540 -180
rect 500 -300 540 -250
rect 620 -180 760 -170
rect 620 -250 630 -180
rect 650 -200 730 -180
rect 750 -200 760 -180
rect 650 -210 760 -200
rect 650 -250 660 -210
rect 620 -260 660 -250
rect -140 -320 60 -300
rect 80 -320 540 -300
rect -140 -340 540 -320
<< labels >>
rlabel metal1 -65 305 -64 306 1 Vdd
rlabel metal1 800 220 820 240 1 vout
rlabel metal1 55 110 55 110 1 VG34
rlabel viali -120 30 -120 30 1 vin2
rlabel metal1 160 -250 160 -250 1 VS12
rlabel metal1 -61 -231 -57 -225 1 vin1
rlabel metal1 170 -330 200 -320 1 Gnd
rlabel metal1 640 -140 650 -130 1 vtail
rlabel metal1 460 60 480 80 1 vinv2
rlabel metal1 322 65 334 75 1 vinv
<< end >>
