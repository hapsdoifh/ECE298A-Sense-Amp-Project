* SPICE3 file created from diff_amp.ext - technology: sky130A

X0 VS12 vin1 VG34 Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X1 vinv VG34 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.84 pd=4 as=0.84 ps=4 w=1.4 l=0.4
X2 voutf Vout2 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.84 pd=4 as=0.84 ps=4 w=1.4 l=0.4
X3 VS12 Vtail Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X4 Vdd VG34 VG34 Vdd sky130_fd_pr__pfet_01v8 ad=0.84 pd=4 as=0.84 ps=4 w=1.4 l=0.4
X5 Vout2 vinv vbase Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X6 voutf Vout2 Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X7 vinv vin2 VS12 Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X8 Vout2 vinv Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.84 pd=4 as=0.84 ps=4 w=1.4 l=0.4
C0 Vdd Gnd 2.30838f
