magic
tech sky130A
timestamp 1763507870
<< nwell >>
rect -100 -20 380 160
<< nmos >>
rect -20 -210 20 -140
rect 260 -210 300 -140
rect 140 -410 180 -340
<< pmos >>
rect -20 0 20 140
rect 260 0 300 140
<< ndiff >>
rect -80 -150 -20 -140
rect -80 -200 -70 -150
rect -50 -200 -20 -150
rect -80 -210 -20 -200
rect 20 -150 80 -140
rect 20 -200 50 -150
rect 70 -200 80 -150
rect 20 -210 80 -200
rect 200 -150 260 -140
rect 200 -200 210 -150
rect 230 -200 260 -150
rect 200 -210 260 -200
rect 300 -150 360 -140
rect 300 -200 330 -150
rect 350 -200 360 -150
rect 300 -210 360 -200
rect 80 -350 140 -340
rect 80 -400 90 -350
rect 110 -400 140 -350
rect 80 -410 140 -400
rect 180 -350 240 -340
rect 180 -400 210 -350
rect 230 -400 240 -350
rect 180 -410 240 -400
<< pdiff >>
rect -80 130 -20 140
rect -80 10 -70 130
rect -50 10 -20 130
rect -80 0 -20 10
rect 20 130 80 140
rect 20 10 50 130
rect 70 10 80 130
rect 200 130 260 140
rect 20 0 80 10
rect 200 10 210 130
rect 230 10 260 130
rect 200 0 260 10
rect 300 130 360 140
rect 300 10 330 130
rect 350 10 360 130
rect 300 0 360 10
<< ndiffc >>
rect -70 -200 -50 -150
rect 50 -200 70 -150
rect 210 -200 230 -150
rect 330 -200 350 -150
rect 90 -400 110 -350
rect 210 -400 230 -350
<< pdiffc >>
rect -70 10 -50 130
rect 50 10 70 130
rect 210 10 230 130
rect 330 10 350 130
<< psubdiff >>
rect -60 -320 20 -300
rect -60 -360 -40 -320
rect 0 -360 20 -320
rect -60 -380 20 -360
<< nsubdiff >>
rect 115 90 165 105
rect 115 70 130 90
rect 150 70 165 90
rect 115 55 165 70
<< psubdiffcont >>
rect -40 -360 0 -320
<< nsubdiffcont >>
rect 130 70 150 90
<< poly >>
rect -20 140 20 170
rect 260 140 300 170
rect -20 -30 20 0
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 260 -30 300 0
rect 260 -50 270 -30
rect 290 -50 300 -30
rect 260 -60 300 -50
rect -20 -100 20 -90
rect -20 -120 -10 -100
rect 10 -120 20 -100
rect -20 -140 20 -120
rect 260 -140 300 -120
rect -20 -230 20 -210
rect 260 -239 300 -210
rect 260 -259 269 -239
rect 290 -259 300 -239
rect 260 -270 300 -259
rect 140 -300 180 -290
rect 140 -320 150 -300
rect 170 -320 180 -300
rect 140 -340 180 -320
rect 140 -430 180 -410
<< polycont >>
rect -10 -50 10 -30
rect 270 -50 290 -30
rect -10 -120 10 -100
rect 269 -259 290 -239
rect 150 -320 170 -300
<< locali >>
rect -80 130 -40 140
rect -80 10 -71 130
rect -50 10 -40 130
rect -80 0 -40 10
rect 40 130 80 140
rect 40 10 50 130
rect 70 10 80 130
rect 200 130 240 140
rect 120 90 160 100
rect 120 70 130 90
rect 150 70 160 90
rect 120 60 160 70
rect 40 0 80 10
rect 200 10 210 130
rect 230 10 240 130
rect 200 0 240 10
rect 320 130 360 140
rect 320 10 330 130
rect 350 10 360 130
rect 320 0 360 10
rect -20 -30 20 -20
rect -20 -50 -10 -30
rect 10 -50 20 -30
rect -20 -60 20 -50
rect 260 -30 300 -20
rect 260 -50 270 -30
rect 290 -50 300 -30
rect 260 -60 300 -50
rect -20 -100 20 -90
rect -20 -120 -10 -100
rect 10 -120 20 -100
rect -20 -130 20 -120
rect -80 -150 -40 -140
rect -80 -200 -70 -150
rect -50 -200 -40 -150
rect -80 -210 -40 -200
rect 40 -150 80 -140
rect 40 -200 50 -150
rect 70 -200 80 -150
rect 40 -210 80 -200
rect 200 -150 240 -140
rect 200 -200 210 -150
rect 230 -200 240 -150
rect 200 -210 240 -200
rect 320 -150 360 -140
rect 320 -200 330 -150
rect 350 -200 360 -150
rect 320 -210 360 -200
rect 260 -239 300 -230
rect 260 -259 269 -239
rect 290 -259 300 -239
rect 260 -270 300 -259
rect 140 -300 180 -290
rect -60 -320 20 -300
rect -60 -360 -40 -320
rect 0 -360 20 -320
rect 140 -320 150 -300
rect 170 -320 180 -300
rect 140 -330 180 -320
rect -60 -380 20 -360
rect 80 -350 120 -340
rect 80 -400 90 -350
rect 110 -400 120 -350
rect 80 -410 120 -400
rect 200 -350 240 -340
rect 200 -400 210 -350
rect 230 -400 240 -350
rect 200 -410 240 -400
<< viali >>
rect -71 10 -70 130
rect -70 10 -50 130
rect 50 10 70 130
rect 130 70 150 90
rect 210 10 230 130
rect 330 10 350 130
rect -10 -50 10 -30
rect 270 -50 290 -30
rect -10 -120 10 -100
rect -70 -200 -50 -150
rect 50 -200 70 -150
rect 210 -200 230 -150
rect 330 -200 350 -150
rect 269 -259 290 -239
rect -40 -360 0 -320
rect 150 -320 170 -300
rect 90 -400 110 -350
rect 210 -400 230 -350
<< metal1 >>
rect -100 230 380 300
rect -80 130 -40 140
rect -80 10 -71 130
rect -50 10 -40 130
rect -80 -20 -40 10
rect 40 130 80 230
rect 40 10 50 130
rect 70 10 80 130
rect 120 90 160 230
rect 120 70 130 90
rect 150 70 160 90
rect 120 60 160 70
rect 200 130 240 230
rect 40 0 80 10
rect 200 10 210 130
rect 230 10 240 130
rect 200 0 240 10
rect 320 130 360 140
rect 320 10 330 130
rect 350 10 360 130
rect -80 -30 300 -20
rect -80 -50 -10 -30
rect 10 -50 270 -30
rect 290 -50 300 -30
rect -80 -60 300 -50
rect -80 -100 20 -90
rect -80 -120 -10 -100
rect 10 -120 20 -100
rect -20 -130 20 -120
rect -80 -150 -40 -140
rect -80 -200 -70 -150
rect -50 -200 -40 -150
rect -80 -230 -40 -200
rect 40 -150 80 -60
rect 40 -200 50 -150
rect 70 -200 80 -150
rect 40 -210 80 -200
rect 200 -150 240 -140
rect 200 -200 210 -150
rect 230 -200 240 -150
rect 200 -230 240 -200
rect 320 -150 360 10
rect 320 -200 330 -150
rect 350 -200 360 -150
rect 320 -210 360 -200
rect -80 -270 240 -230
rect 260 -239 360 -230
rect 260 -259 269 -239
rect 290 -259 360 -239
rect 260 -270 360 -259
rect 80 -300 180 -290
rect -60 -320 20 -300
rect 80 -320 150 -300
rect 170 -320 180 -300
rect -60 -360 -40 -320
rect 0 -360 20 -320
rect 140 -330 180 -320
rect -60 -440 20 -360
rect 80 -350 120 -340
rect 80 -400 90 -350
rect 110 -400 120 -350
rect 80 -440 120 -400
rect 200 -350 240 -270
rect 200 -400 210 -350
rect 230 -400 240 -350
rect 200 -410 240 -400
rect -100 -441 380 -440
rect -101 -510 380 -441
<< labels >>
rlabel metal1 -65 265 -64 266 1 Vdd
rlabel metal1 55 -40 55 -40 1 VG34
rlabel metal1 340 -250 340 -250 1 Vin2
rlabel metal1 -65 -110 -65 -110 1 Vin1
rlabel metal1 94 -307 95 -306 1 Vtail
rlabel metal1 -3 -252 -3 -252 1 VD12
rlabel metal1 341 -76 341 -76 1 Vout
rlabel metal1 90 -480 93 -477 1 Gnd
<< end >>
