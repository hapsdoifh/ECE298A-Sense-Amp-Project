* SPICE3 file created from diff_amp.ext - technology: sky130A

X0 vinv VG34 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.72 pd=3.6 as=0.72 ps=3.6 w=1.2 l=0.4
X1 VS12 vin1 VG34 Gnd sky130_fd_pr__nfet_01v8 ad=0.96 pd=4.4 as=0.96 ps=4.4 w=1.6 l=0.4
X2 vinv2 vinv Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.72 pd=3.6 as=0.72 ps=3.6 w=1.2 l=0.4
X3 vout vinv2 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=5.4 as=1.26 ps=5.4 w=2.1 l=0.4
X4 Vdd VG34 VG34 Vdd sky130_fd_pr__pfet_01v8 ad=0.72 pd=3.6 as=0.72 ps=3.6 w=1.2 l=0.4
X5 vinv vin2 VS12 Gnd sky130_fd_pr__nfet_01v8 ad=0.96 pd=4.4 as=0.96 ps=4.4 w=1.6 l=0.4
X6 vout vinv2 Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.72 pd=3.6 as=0.72 ps=3.6 w=1.2 l=0.4
X7 vtail vtail Gnd Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
X8 vinv2 vinv Vdd Vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=5.4 as=1.26 ps=5.4 w=2.1 l=0.4
X9 Vdd vtail Gnd sky130_fd_pr__res_xhigh_po w=0.4 l=1.06
X10 Gnd vtail VS12 Gnd sky130_fd_pr__nfet_01v8 ad=0.42 pd=2.6 as=0.42 ps=2.6 w=0.7 l=0.4
C0 Vdd Gnd 3.30401f 
