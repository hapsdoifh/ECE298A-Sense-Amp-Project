magic
tech sky130A
timestamp 1764711567
<< nwell >>
rect 40 230 150 310
rect -100 130 680 230
rect 270 70 680 130
<< nmos >>
rect 370 -40 410 10
rect 560 -40 600 10
rect -20 -270 20 -60
rect 170 -270 210 -60
rect 370 -340 410 -190
rect 560 -340 600 -190
<< pmos >>
rect -20 150 20 210
rect 170 150 210 210
rect 370 90 410 210
rect 560 90 600 210
<< ndiff >>
rect 310 0 370 10
rect 310 -30 320 0
rect 340 -30 370 0
rect 310 -40 370 -30
rect 410 0 470 10
rect 410 -30 440 0
rect 460 -30 470 0
rect 410 -40 470 -30
rect 500 0 560 10
rect 500 -30 510 0
rect 530 -30 560 0
rect 500 -40 560 -30
rect 600 0 660 10
rect 600 -30 630 0
rect 650 -30 660 0
rect 600 -40 660 -30
rect -80 -70 -20 -60
rect -80 -260 -70 -70
rect -50 -260 -20 -70
rect -80 -270 -20 -260
rect 20 -70 80 -60
rect 20 -260 50 -70
rect 70 -260 80 -70
rect 20 -270 80 -260
rect 110 -70 170 -60
rect 110 -260 120 -70
rect 140 -260 170 -70
rect 110 -270 170 -260
rect 210 -70 270 -60
rect 210 -260 240 -70
rect 260 -260 270 -70
rect 210 -270 270 -260
rect 310 -200 370 -190
rect 310 -330 320 -200
rect 340 -330 370 -200
rect 310 -340 370 -330
rect 410 -200 470 -190
rect 410 -330 440 -200
rect 460 -330 470 -200
rect 410 -340 470 -330
rect 500 -200 560 -190
rect 500 -330 510 -200
rect 530 -330 560 -200
rect 500 -340 560 -330
rect 600 -200 660 -190
rect 600 -330 630 -200
rect 650 -330 660 -200
rect 600 -340 660 -330
<< pdiff >>
rect -80 200 -20 210
rect -80 160 -70 200
rect -50 160 -20 200
rect -80 150 -20 160
rect 20 200 80 210
rect 20 160 50 200
rect 70 160 80 200
rect 20 150 80 160
rect 110 200 170 210
rect 110 160 120 200
rect 140 160 170 200
rect 110 150 170 160
rect 210 200 270 210
rect 210 160 240 200
rect 260 160 270 200
rect 210 150 270 160
rect 310 200 370 210
rect 310 100 320 200
rect 340 100 370 200
rect 310 90 370 100
rect 410 200 470 210
rect 410 100 440 200
rect 460 100 470 200
rect 410 90 470 100
rect 500 200 560 210
rect 500 100 510 200
rect 530 100 560 200
rect 500 90 560 100
rect 600 200 660 210
rect 600 100 630 200
rect 650 100 660 200
rect 600 90 660 100
<< ndiffc >>
rect 320 -30 340 0
rect 440 -30 460 0
rect 510 -30 530 0
rect 630 -30 650 0
rect -70 -260 -50 -70
rect 50 -260 70 -70
rect 120 -260 140 -70
rect 240 -260 260 -70
rect 320 -330 340 -200
rect 440 -330 460 -200
rect 510 -330 530 -200
rect 630 -330 650 -200
<< pdiffc >>
rect -70 160 -50 200
rect 50 160 70 200
rect 120 160 140 200
rect 240 160 260 200
rect 320 100 340 200
rect 440 100 460 200
rect 510 100 530 200
rect 630 100 650 200
<< psubdiff >>
rect -100 -380 -40 -360
rect -100 -400 -80 -380
rect -60 -400 -40 -380
rect -100 -420 -40 -400
<< nsubdiff >>
rect 75 275 115 290
rect 75 255 85 275
rect 105 255 115 275
rect 75 240 115 255
<< psubdiffcont >>
rect -80 -400 -60 -380
<< nsubdiffcont >>
rect 85 255 105 275
<< poly >>
rect -20 210 20 240
rect 170 210 210 240
rect 370 210 410 240
rect 560 210 600 240
rect -20 120 20 150
rect -20 100 -10 120
rect 10 100 20 120
rect -20 90 20 100
rect 170 120 210 150
rect 170 100 180 120
rect 200 100 210 120
rect 170 90 210 100
rect 370 60 410 90
rect 370 40 380 60
rect 400 40 410 60
rect 370 10 410 40
rect 560 60 600 90
rect 560 40 570 60
rect 590 40 600 60
rect 560 10 600 40
rect 170 -10 210 0
rect 170 -30 180 -10
rect 200 -30 210 -10
rect -20 -60 20 -40
rect 170 -60 210 -30
rect 370 -60 410 -40
rect 560 -60 600 -40
rect 370 -140 410 -130
rect 370 -160 380 -140
rect 400 -160 410 -140
rect 370 -190 410 -160
rect 560 -140 600 -130
rect 560 -160 570 -140
rect 590 -160 600 -140
rect 560 -190 600 -160
rect -20 -299 20 -270
rect 170 -290 210 -270
rect -20 -319 -11 -299
rect 10 -319 20 -299
rect -20 -330 20 -319
rect 370 -360 410 -340
rect 560 -360 600 -340
<< polycont >>
rect -10 100 10 120
rect 180 100 200 120
rect 380 40 400 60
rect 570 40 590 60
rect 180 -30 200 -10
rect 380 -160 400 -140
rect 570 -160 590 -140
rect -11 -319 10 -299
<< xpolycontact >>
rect 720 70 760 310
rect 720 -210 760 30
<< xpolyres >>
rect 720 30 760 70
<< locali >>
rect 75 275 115 285
rect 75 255 85 275
rect 105 255 115 275
rect 75 245 115 255
rect -80 200 -40 210
rect -80 160 -70 200
rect -50 160 -40 200
rect -80 150 -40 160
rect 40 200 80 210
rect 40 160 50 200
rect 70 160 80 200
rect 40 150 80 160
rect 110 200 150 210
rect 110 160 120 200
rect 140 160 150 200
rect 110 150 150 160
rect 230 200 270 210
rect 230 160 240 200
rect 260 160 270 200
rect 230 150 270 160
rect 310 200 350 210
rect -20 120 20 130
rect -20 100 -10 120
rect 10 100 20 120
rect -20 90 20 100
rect 170 120 210 130
rect 170 100 180 120
rect 200 100 210 120
rect 170 90 210 100
rect 310 100 320 200
rect 340 100 350 200
rect 310 90 350 100
rect 430 200 470 210
rect 430 100 440 200
rect 460 100 470 200
rect 430 90 470 100
rect 500 200 540 210
rect 500 100 510 200
rect 530 100 540 200
rect 500 90 540 100
rect 620 200 660 210
rect 620 100 630 200
rect 650 100 660 200
rect 620 90 660 100
rect 370 60 410 70
rect 370 40 380 60
rect 400 40 410 60
rect 370 30 410 40
rect 560 60 600 70
rect 560 40 570 60
rect 590 40 600 60
rect 560 30 600 40
rect 310 0 350 10
rect -140 -10 20 0
rect -140 -30 -130 -10
rect -110 -30 -10 -10
rect 10 -30 20 -10
rect -140 -40 20 -30
rect 170 -10 210 0
rect 170 -30 180 -10
rect 200 -30 210 -10
rect 170 -40 210 -30
rect 310 -30 320 0
rect 340 -30 350 0
rect 310 -40 350 -30
rect 430 0 470 10
rect 430 -30 440 0
rect 460 -30 470 0
rect 430 -40 470 -30
rect 500 0 540 10
rect 500 -30 510 0
rect 530 -30 540 0
rect 500 -40 540 -30
rect 620 0 660 10
rect 620 -30 630 0
rect 650 -30 660 0
rect 620 -40 660 -30
rect -80 -70 -40 -60
rect -80 -260 -70 -70
rect -50 -260 -40 -70
rect -80 -270 -40 -260
rect 40 -70 80 -60
rect 40 -260 50 -70
rect 70 -260 80 -70
rect 40 -270 80 -260
rect 110 -70 150 -60
rect 110 -260 120 -70
rect 140 -260 150 -70
rect 110 -270 150 -260
rect 230 -70 270 -60
rect 230 -260 240 -70
rect 260 -260 270 -70
rect 500 -80 540 -70
rect 500 -100 510 -80
rect 530 -100 540 -80
rect 370 -140 410 -130
rect 370 -160 380 -140
rect 400 -160 410 -140
rect 370 -170 410 -160
rect 230 -270 270 -260
rect 310 -200 350 -190
rect -20 -299 20 -290
rect -20 -319 -11 -299
rect 10 -319 20 -299
rect -20 -330 20 -319
rect 310 -330 320 -200
rect 340 -330 350 -200
rect 310 -340 350 -330
rect 430 -200 470 -190
rect 430 -330 440 -200
rect 460 -330 470 -200
rect 430 -340 470 -330
rect 500 -200 540 -100
rect 560 -140 600 -130
rect 560 -160 570 -140
rect 590 -160 600 -140
rect 560 -170 600 -160
rect 500 -330 510 -200
rect 530 -330 540 -200
rect 500 -340 540 -330
rect 620 -200 660 -190
rect 620 -330 630 -200
rect 650 -330 660 -200
rect 620 -340 660 -330
rect -100 -380 -40 -360
rect -100 -400 -80 -380
rect -60 -400 -40 -380
rect -100 -420 -40 -400
<< viali >>
rect 85 255 105 275
rect 730 280 750 300
rect -70 160 -50 200
rect 50 160 70 200
rect 120 160 140 200
rect 240 160 260 200
rect -10 100 10 120
rect 180 100 200 120
rect 320 100 340 200
rect 440 100 460 200
rect 510 100 530 200
rect 630 100 650 200
rect 380 40 400 60
rect 570 40 590 60
rect -130 -30 -110 -10
rect -10 -30 10 -10
rect 180 -30 200 -10
rect 320 -30 340 0
rect 440 -30 460 0
rect 510 -30 530 0
rect 630 -30 650 0
rect -70 -260 -50 -70
rect 50 -260 70 -70
rect 120 -260 140 -70
rect 240 -260 260 -70
rect 510 -100 530 -80
rect 380 -160 400 -140
rect -11 -319 10 -299
rect 320 -330 340 -200
rect 440 -330 460 -200
rect 570 -160 590 -140
rect 510 -330 530 -200
rect 630 -330 650 -200
rect 730 -200 750 -180
rect -80 -400 -60 -380
<< metal1 >>
rect -140 300 760 310
rect -140 280 730 300
rect 750 280 760 300
rect -140 275 760 280
rect -140 270 85 275
rect 40 255 85 270
rect 105 270 760 275
rect 105 255 150 270
rect 40 230 150 255
rect -80 200 -40 210
rect -80 160 -70 200
rect -50 160 -40 200
rect -80 130 -40 160
rect 40 200 80 230
rect 40 160 50 200
rect 70 160 80 200
rect 40 150 80 160
rect 110 200 150 230
rect 110 160 120 200
rect 140 160 150 200
rect 110 150 150 160
rect 230 200 270 210
rect 230 160 240 200
rect 260 160 270 200
rect -80 120 210 130
rect -80 100 -10 120
rect 10 100 180 120
rect 200 100 210 120
rect -80 90 210 100
rect -140 -10 -100 0
rect -140 -30 -130 -10
rect -110 -30 -100 -10
rect -140 -40 -100 -30
rect -80 -70 -40 90
rect 230 70 270 160
rect 310 200 350 270
rect 310 100 320 200
rect 340 100 350 200
rect 310 90 350 100
rect 430 200 470 210
rect 430 100 440 200
rect 460 100 470 200
rect 230 60 410 70
rect 230 40 380 60
rect 400 40 410 60
rect 230 30 410 40
rect 430 69 470 100
rect 500 200 540 270
rect 500 100 510 200
rect 530 100 540 200
rect 500 90 540 100
rect 620 210 830 250
rect 620 200 660 210
rect 620 100 630 200
rect 650 100 660 200
rect 500 69 600 70
rect 430 60 600 69
rect 430 40 570 60
rect 590 40 600 60
rect 430 30 600 40
rect -20 -10 210 0
rect -20 -30 -10 -10
rect 10 -30 180 -10
rect 200 -30 210 -10
rect -20 -40 210 -30
rect -80 -260 -70 -70
rect -50 -260 -40 -70
rect -80 -270 -40 -260
rect 40 -70 80 -60
rect 40 -260 50 -70
rect 70 -250 80 -70
rect 110 -70 150 -60
rect 110 -250 120 -70
rect 70 -260 120 -250
rect 140 -260 150 -70
rect 40 -270 150 -260
rect 230 -70 270 30
rect 230 -260 240 -70
rect 260 -260 270 -70
rect 310 0 350 10
rect 310 -30 320 0
rect 340 -30 350 0
rect 310 -70 350 -30
rect 430 0 470 30
rect 430 -30 440 0
rect 460 -30 470 0
rect 430 -40 470 -30
rect 500 0 540 10
rect 500 -30 510 0
rect 530 -30 540 0
rect 500 -70 540 -30
rect 620 0 660 100
rect 620 -30 630 0
rect 650 -30 660 0
rect 620 -40 660 -30
rect 310 -80 540 -70
rect 310 -100 510 -80
rect 530 -100 540 -80
rect 310 -110 540 -100
rect 370 -140 660 -130
rect 370 -160 380 -140
rect 400 -160 570 -140
rect 590 -160 660 -140
rect 370 -170 660 -160
rect 620 -180 760 -170
rect 230 -270 270 -260
rect 310 -200 350 -190
rect -140 -299 20 -290
rect -140 -319 -11 -299
rect 10 -319 20 -299
rect -140 -330 20 -319
rect 110 -300 150 -270
rect 310 -300 320 -200
rect 110 -330 320 -300
rect 340 -330 350 -200
rect 110 -340 350 -330
rect 430 -200 470 -190
rect 430 -330 440 -200
rect 460 -330 470 -200
rect -100 -380 -40 -360
rect 430 -380 470 -330
rect 500 -200 540 -190
rect 500 -330 510 -200
rect 530 -330 540 -200
rect 500 -380 540 -330
rect 620 -200 730 -180
rect 750 -200 760 -180
rect 620 -330 630 -200
rect 650 -210 760 -200
rect 650 -330 660 -210
rect 620 -340 660 -330
rect -140 -400 -80 -380
rect -60 -400 540 -380
rect -140 -420 540 -400
<< labels >>
rlabel metal1 -65 305 -64 306 1 Vdd
rlabel metal1 640 -160 650 -150 1 vtail
rlabel metal1 460 40 480 60 1 vinv2
rlabel metal1 322 45 334 55 1 vinv
rlabel metal1 800 220 820 240 1 vout
rlabel viali -120 -20 -120 -20 1 vin2
rlabel metal1 170 -410 200 -400 1 Gnd
rlabel metal1 160 -330 160 -330 1 VS12
rlabel metal1 -61 -311 -57 -305 1 vin1
rlabel metal1 55 110 55 110 1 VG34
<< end >>
