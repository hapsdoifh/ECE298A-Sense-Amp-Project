magic
tech sky130A
timestamp 1764652427
<< nwell >>
rect 40 230 150 310
rect -100 30 690 230
rect 270 -20 690 30
<< nmos >>
rect -20 -220 20 -100
rect 170 -220 210 -100
rect 370 -130 410 -80
rect 570 -130 610 -80
rect 100 -440 140 -370
rect 290 -440 330 -370
<< pmos >>
rect -20 50 20 210
rect 170 50 210 210
rect 370 0 410 210
rect 570 0 610 210
<< ndiff >>
rect 310 -90 370 -80
rect -80 -110 -20 -100
rect -80 -210 -70 -110
rect -50 -210 -20 -110
rect -80 -220 -20 -210
rect 20 -110 80 -100
rect 20 -210 50 -110
rect 70 -210 80 -110
rect 20 -220 80 -210
rect 110 -110 170 -100
rect 110 -210 120 -110
rect 140 -210 170 -110
rect 110 -220 170 -210
rect 210 -110 270 -100
rect 210 -210 240 -110
rect 260 -210 270 -110
rect 310 -120 320 -90
rect 340 -120 370 -90
rect 310 -130 370 -120
rect 410 -90 470 -80
rect 410 -120 440 -90
rect 460 -120 470 -90
rect 410 -130 470 -120
rect 510 -90 570 -80
rect 510 -120 520 -90
rect 540 -120 570 -90
rect 510 -130 570 -120
rect 610 -90 670 -80
rect 610 -120 640 -90
rect 660 -120 670 -90
rect 610 -130 670 -120
rect 210 -220 270 -210
rect 40 -380 100 -370
rect 40 -430 50 -380
rect 70 -430 100 -380
rect 40 -440 100 -430
rect 140 -380 200 -370
rect 140 -430 170 -380
rect 190 -430 200 -380
rect 140 -440 200 -430
rect 230 -380 290 -370
rect 230 -430 240 -380
rect 260 -430 290 -380
rect 230 -440 290 -430
rect 330 -380 390 -370
rect 330 -430 360 -380
rect 380 -430 390 -380
rect 330 -440 390 -430
<< pdiff >>
rect -80 200 -20 210
rect -80 60 -70 200
rect -50 60 -20 200
rect -80 50 -20 60
rect 20 200 80 210
rect 20 60 50 200
rect 70 60 80 200
rect 20 50 80 60
rect 110 200 170 210
rect 110 60 120 200
rect 140 60 170 200
rect 110 50 170 60
rect 210 200 270 210
rect 210 60 240 200
rect 260 60 270 200
rect 210 50 270 60
rect 310 200 370 210
rect 310 10 320 200
rect 340 10 370 200
rect 310 0 370 10
rect 410 200 470 210
rect 410 10 440 200
rect 460 10 470 200
rect 410 0 470 10
rect 510 200 570 210
rect 510 10 520 200
rect 540 10 570 200
rect 510 0 570 10
rect 610 200 670 210
rect 610 10 640 200
rect 660 10 670 200
rect 610 0 670 10
<< ndiffc >>
rect -70 -210 -50 -110
rect 50 -210 70 -110
rect 120 -210 140 -110
rect 240 -210 260 -110
rect 320 -120 340 -90
rect 440 -120 460 -90
rect 520 -120 540 -90
rect 640 -120 660 -90
rect 50 -430 70 -380
rect 170 -430 190 -380
rect 240 -430 260 -380
rect 360 -430 380 -380
<< pdiffc >>
rect -70 60 -50 200
rect 50 60 70 200
rect 120 60 140 200
rect 240 60 260 200
rect 320 10 340 200
rect 440 10 460 200
rect 520 10 540 200
rect 640 10 660 200
<< psubdiff >>
rect -100 -400 -40 -380
rect -100 -420 -80 -400
rect -60 -420 -40 -400
rect -100 -440 -40 -420
<< nsubdiff >>
rect 75 275 115 290
rect 75 255 85 275
rect 105 255 115 275
rect 75 240 115 255
<< psubdiffcont >>
rect -80 -420 -60 -400
<< nsubdiffcont >>
rect 85 255 105 275
<< poly >>
rect -20 210 20 240
rect 170 210 210 240
rect 370 210 410 240
rect 570 210 610 240
rect -20 20 20 50
rect -20 0 -10 20
rect 10 0 20 20
rect -20 -10 20 0
rect 170 20 210 50
rect 170 0 180 20
rect 200 0 210 20
rect 170 -10 210 0
rect 370 -30 410 0
rect 170 -50 210 -40
rect 170 -70 180 -50
rect 200 -70 210 -50
rect -20 -100 20 -80
rect 170 -100 210 -70
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -80 410 -50
rect 570 -30 610 0
rect 570 -50 580 -30
rect 600 -50 610 -30
rect 570 -80 610 -50
rect 370 -150 410 -130
rect 570 -150 610 -130
rect -20 -249 20 -220
rect 170 -240 210 -220
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 100 -320 140 -310
rect 100 -340 110 -320
rect 130 -340 140 -320
rect 100 -370 140 -340
rect 290 -320 330 -310
rect 290 -340 300 -320
rect 320 -340 330 -320
rect 290 -370 330 -340
rect 100 -460 140 -440
rect 290 -460 330 -440
<< polycont >>
rect -10 0 10 20
rect 180 0 200 20
rect 180 -70 200 -50
rect 380 -50 400 -30
rect 580 -50 600 -30
rect -11 -269 10 -249
rect 110 -340 130 -320
rect 300 -340 320 -320
<< xpolycontact >>
rect 730 -310 770 30
rect 450 -350 670 -310
<< xpolyres >>
rect 670 -350 770 -310
<< locali >>
rect 730 300 770 310
rect 75 275 115 285
rect 75 255 85 275
rect 105 255 115 275
rect 75 245 115 255
rect 730 280 740 300
rect 760 280 770 300
rect -80 200 -40 210
rect -80 60 -70 200
rect -50 60 -40 200
rect -80 50 -40 60
rect 40 200 80 210
rect 40 60 50 200
rect 70 60 80 200
rect 40 50 80 60
rect 110 200 150 210
rect 110 60 120 200
rect 140 60 150 200
rect 110 50 150 60
rect 230 200 270 210
rect 230 60 240 200
rect 260 60 270 200
rect 230 50 270 60
rect 310 200 350 210
rect -20 20 20 30
rect -20 0 -10 20
rect 10 0 20 20
rect -20 -10 20 0
rect 170 20 210 30
rect 170 0 180 20
rect 200 0 210 20
rect 310 10 320 200
rect 340 10 350 200
rect 310 0 350 10
rect 430 200 470 210
rect 430 10 440 200
rect 460 10 470 200
rect 430 0 470 10
rect 510 200 550 210
rect 510 10 520 200
rect 540 10 550 200
rect 510 0 550 10
rect 630 200 670 210
rect 630 10 640 200
rect 660 10 670 200
rect 730 180 770 280
rect 730 160 740 180
rect 760 160 770 180
rect 730 150 770 160
rect 630 0 670 10
rect 170 -10 210 0
rect 370 -30 410 -20
rect -140 -50 20 -40
rect -140 -70 -130 -50
rect -110 -70 -10 -50
rect 10 -70 20 -50
rect -140 -80 20 -70
rect 170 -50 210 -40
rect 170 -70 180 -50
rect 200 -70 210 -50
rect 370 -50 380 -30
rect 400 -50 410 -30
rect 370 -60 410 -50
rect 570 -30 610 -20
rect 570 -50 580 -30
rect 600 -50 610 -30
rect 570 -60 610 -50
rect 170 -80 210 -70
rect 310 -90 350 -80
rect -80 -110 -40 -100
rect -80 -210 -70 -110
rect -50 -210 -40 -110
rect -80 -220 -40 -210
rect 40 -110 80 -100
rect 40 -210 50 -110
rect 70 -210 80 -110
rect 40 -220 80 -210
rect 110 -110 150 -100
rect 110 -210 120 -110
rect 140 -210 150 -110
rect 110 -220 150 -210
rect 230 -110 270 -100
rect 230 -210 240 -110
rect 260 -210 270 -110
rect 310 -120 320 -90
rect 340 -120 350 -90
rect 310 -130 350 -120
rect 430 -90 470 -80
rect 430 -120 440 -90
rect 460 -120 470 -90
rect 430 -130 470 -120
rect 510 -90 550 -80
rect 510 -120 520 -90
rect 540 -120 550 -90
rect 510 -130 550 -120
rect 630 -90 670 -80
rect 630 -120 640 -90
rect 660 -120 670 -90
rect 630 -130 670 -120
rect 230 -220 270 -210
rect -20 -249 20 -240
rect -20 -269 -11 -249
rect 10 -269 20 -249
rect -20 -280 20 -269
rect 100 -320 140 -310
rect 100 -340 110 -320
rect 130 -340 140 -320
rect 100 -350 140 -340
rect 290 -320 330 -310
rect 290 -340 300 -320
rect 320 -340 330 -320
rect 290 -350 330 -340
rect 40 -380 80 -370
rect -100 -400 -40 -380
rect -100 -420 -80 -400
rect -60 -420 -40 -400
rect -100 -440 -40 -420
rect 40 -430 50 -380
rect 70 -430 80 -380
rect 40 -440 80 -430
rect 160 -380 200 -370
rect 160 -430 170 -380
rect 190 -430 200 -380
rect 160 -440 200 -430
rect 230 -380 270 -370
rect 230 -430 240 -380
rect 260 -430 270 -380
rect 230 -440 270 -430
rect 350 -380 390 -370
rect 350 -430 360 -380
rect 380 -430 390 -380
rect 350 -440 390 -430
<< viali >>
rect 85 255 105 275
rect 740 280 760 300
rect -70 60 -50 200
rect 50 60 70 200
rect 120 60 140 200
rect 240 60 260 200
rect -10 0 10 20
rect 180 0 200 20
rect 320 10 340 200
rect 440 10 460 200
rect 520 10 540 200
rect 640 10 660 200
rect 740 160 760 180
rect 740 0 760 20
rect -130 -70 -110 -50
rect -10 -70 10 -50
rect 180 -70 200 -50
rect 380 -50 400 -30
rect 580 -50 600 -30
rect -70 -210 -50 -110
rect 50 -210 70 -110
rect 120 -210 140 -110
rect 240 -210 260 -110
rect 320 -120 340 -90
rect 440 -120 460 -90
rect 520 -120 540 -90
rect 640 -120 660 -90
rect -11 -269 10 -249
rect 110 -340 130 -320
rect 300 -340 320 -320
rect 460 -340 480 -320
rect -80 -420 -60 -400
rect 50 -430 70 -380
rect 170 -430 190 -380
rect 240 -430 260 -380
rect 360 -430 380 -380
<< metal1 >>
rect -140 300 770 310
rect -140 280 740 300
rect 760 280 770 300
rect -140 275 770 280
rect -140 270 85 275
rect 40 255 85 270
rect 105 270 770 275
rect 105 255 150 270
rect 40 230 150 255
rect -80 200 -40 210
rect -80 60 -70 200
rect -50 60 -40 200
rect -80 30 -40 60
rect 40 200 80 230
rect 40 60 50 200
rect 70 60 80 200
rect 40 50 80 60
rect 110 200 150 230
rect 110 60 120 200
rect 140 60 150 200
rect 110 50 150 60
rect 230 200 270 210
rect 230 60 240 200
rect 260 60 270 200
rect -80 20 210 30
rect -80 0 -10 20
rect 10 0 180 20
rect 200 0 210 20
rect -80 -10 210 0
rect -140 -50 -100 -40
rect -140 -70 -130 -50
rect -110 -70 -100 -50
rect -140 -80 -100 -70
rect -80 -110 -40 -10
rect 230 -20 270 60
rect 310 200 350 270
rect 310 10 320 200
rect 340 10 350 200
rect 310 0 350 10
rect 430 200 470 210
rect 430 10 440 200
rect 460 10 470 200
rect 230 -30 410 -20
rect -20 -50 210 -40
rect -20 -70 -10 -50
rect 10 -70 180 -50
rect 200 -70 210 -50
rect -20 -80 210 -70
rect 230 -50 380 -30
rect 400 -50 410 -30
rect 230 -60 410 -50
rect 430 -21 470 10
rect 510 200 550 270
rect 510 10 520 200
rect 540 10 550 200
rect 510 0 550 10
rect 630 210 840 250
rect 630 200 670 210
rect 630 10 640 200
rect 660 10 670 200
rect 510 -21 610 -20
rect 430 -30 610 -21
rect 430 -50 580 -30
rect 600 -50 610 -30
rect 430 -60 610 -50
rect -80 -210 -70 -110
rect -50 -210 -40 -110
rect -80 -220 -40 -210
rect 40 -110 80 -100
rect 40 -210 50 -110
rect 70 -210 80 -110
rect 110 -110 150 -100
rect 110 -210 120 -110
rect 140 -210 150 -110
rect -140 -249 20 -240
rect -140 -269 -11 -249
rect 10 -269 20 -249
rect -140 -280 20 -269
rect 40 -260 150 -210
rect 230 -110 270 -60
rect 230 -210 240 -110
rect 260 -210 270 -110
rect 230 -220 270 -210
rect 310 -90 350 -80
rect 310 -120 320 -90
rect 340 -120 350 -90
rect 310 -250 350 -120
rect 430 -90 470 -60
rect 430 -120 440 -90
rect 460 -120 470 -90
rect 430 -130 470 -120
rect 510 -90 550 -80
rect 510 -120 520 -90
rect 540 -120 550 -90
rect 510 -190 550 -120
rect 630 -90 670 10
rect 730 180 770 190
rect 730 160 740 180
rect 760 160 770 180
rect 730 20 770 160
rect 730 0 740 20
rect 760 0 770 20
rect 730 -10 770 0
rect 630 -120 640 -90
rect 660 -120 670 -90
rect 630 -130 670 -120
rect 510 -230 670 -190
rect 40 -380 80 -260
rect 310 -290 610 -250
rect 100 -320 490 -310
rect 100 -340 110 -320
rect 130 -340 300 -320
rect 320 -340 460 -320
rect 480 -340 490 -320
rect 100 -350 490 -340
rect -100 -400 -40 -380
rect -100 -420 -80 -400
rect -60 -420 -40 -400
rect -100 -480 -40 -420
rect 40 -430 50 -380
rect 70 -430 80 -380
rect 40 -440 80 -430
rect 160 -380 200 -370
rect 160 -430 170 -380
rect 190 -430 200 -380
rect 160 -480 200 -430
rect 230 -380 270 -370
rect 230 -430 240 -380
rect 260 -430 270 -380
rect 230 -480 270 -430
rect 350 -380 390 -350
rect 350 -430 360 -380
rect 380 -430 390 -380
rect 350 -440 390 -430
rect 570 -370 610 -290
rect 630 -370 670 -230
rect 570 -480 670 -370
rect -140 -520 670 -480
<< labels >>
rlabel metal1 -65 305 -64 306 1 Vdd
rlabel metal1 322 -45 334 -35 1 vinv
rlabel metal1 460 -50 480 -30 1 vinv2
rlabel metal1 90 -230 90 -230 1 VS12
rlabel metal1 -61 -261 -57 -255 1 vin1
rlabel metal1 55 10 55 10 1 VG34
rlabel viali -120 -60 -120 -60 1 vin2
rlabel metal1 810 220 830 240 1 vout
rlabel metal1 170 -510 200 -500 1 Gnd
<< end >>
